// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire net220;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net221;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net222;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net258;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net278;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net279;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net280;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net281;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net282;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net283;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire \mod.clk ;
 wire \mod.des.des_counter[0] ;
 wire \mod.des.des_counter[1] ;
 wire \mod.des.des_counter[2] ;
 wire \mod.des.des_dout[0] ;
 wire \mod.des.des_dout[10] ;
 wire \mod.des.des_dout[11] ;
 wire \mod.des.des_dout[12] ;
 wire \mod.des.des_dout[13] ;
 wire \mod.des.des_dout[14] ;
 wire \mod.des.des_dout[15] ;
 wire \mod.des.des_dout[16] ;
 wire \mod.des.des_dout[17] ;
 wire \mod.des.des_dout[18] ;
 wire \mod.des.des_dout[19] ;
 wire \mod.des.des_dout[1] ;
 wire \mod.des.des_dout[20] ;
 wire \mod.des.des_dout[21] ;
 wire \mod.des.des_dout[22] ;
 wire \mod.des.des_dout[23] ;
 wire \mod.des.des_dout[24] ;
 wire \mod.des.des_dout[25] ;
 wire \mod.des.des_dout[26] ;
 wire \mod.des.des_dout[27] ;
 wire \mod.des.des_dout[28] ;
 wire \mod.des.des_dout[29] ;
 wire \mod.des.des_dout[2] ;
 wire \mod.des.des_dout[30] ;
 wire \mod.des.des_dout[31] ;
 wire \mod.des.des_dout[32] ;
 wire \mod.des.des_dout[33] ;
 wire \mod.des.des_dout[34] ;
 wire \mod.des.des_dout[35] ;
 wire \mod.des.des_dout[36] ;
 wire \mod.des.des_dout[3] ;
 wire \mod.des.des_dout[4] ;
 wire \mod.des.des_dout[5] ;
 wire \mod.des.des_dout[6] ;
 wire \mod.des.des_dout[7] ;
 wire \mod.des.des_dout[8] ;
 wire \mod.des.des_dout[9] ;
 wire \mod.funct3[0] ;
 wire \mod.funct3[1] ;
 wire \mod.funct3[2] ;
 wire \mod.funct7[0] ;
 wire \mod.funct7[1] ;
 wire \mod.funct7[2] ;
 wire \mod.ins_ldr_3 ;
 wire \mod.instr[0] ;
 wire \mod.instr[10] ;
 wire \mod.instr[11] ;
 wire \mod.instr[12] ;
 wire \mod.instr[13] ;
 wire \mod.instr[14] ;
 wire \mod.instr[15] ;
 wire \mod.instr[16] ;
 wire \mod.instr[17] ;
 wire \mod.instr[18] ;
 wire \mod.instr[19] ;
 wire \mod.instr[1] ;
 wire \mod.instr[20] ;
 wire \mod.instr[2] ;
 wire \mod.instr[3] ;
 wire \mod.instr[4] ;
 wire \mod.instr[5] ;
 wire \mod.instr[6] ;
 wire \mod.instr[7] ;
 wire \mod.instr[8] ;
 wire \mod.instr[9] ;
 wire \mod.instr_2[0] ;
 wire \mod.instr_2[10] ;
 wire \mod.instr_2[11] ;
 wire \mod.instr_2[12] ;
 wire \mod.instr_2[13] ;
 wire \mod.instr_2[14] ;
 wire \mod.instr_2[15] ;
 wire \mod.instr_2[16] ;
 wire \mod.instr_2[17] ;
 wire \mod.instr_2[1] ;
 wire \mod.instr_2[2] ;
 wire \mod.instr_2[3] ;
 wire \mod.instr_2[4] ;
 wire \mod.instr_2[5] ;
 wire \mod.instr_2[6] ;
 wire \mod.ldr_hzd[0] ;
 wire \mod.ldr_hzd[10] ;
 wire \mod.ldr_hzd[11] ;
 wire \mod.ldr_hzd[12] ;
 wire \mod.ldr_hzd[13] ;
 wire \mod.ldr_hzd[14] ;
 wire \mod.ldr_hzd[15] ;
 wire \mod.ldr_hzd[1] ;
 wire \mod.ldr_hzd[2] ;
 wire \mod.ldr_hzd[3] ;
 wire \mod.ldr_hzd[4] ;
 wire \mod.ldr_hzd[5] ;
 wire \mod.ldr_hzd[6] ;
 wire \mod.ldr_hzd[7] ;
 wire \mod.ldr_hzd[8] ;
 wire \mod.ldr_hzd[9] ;
 wire \mod.pc0[0] ;
 wire \mod.pc0[10] ;
 wire \mod.pc0[11] ;
 wire \mod.pc0[12] ;
 wire \mod.pc0[13] ;
 wire \mod.pc0[1] ;
 wire \mod.pc0[2] ;
 wire \mod.pc0[3] ;
 wire \mod.pc0[4] ;
 wire \mod.pc0[5] ;
 wire \mod.pc0[6] ;
 wire \mod.pc0[7] ;
 wire \mod.pc0[8] ;
 wire \mod.pc0[9] ;
 wire \mod.pc[0] ;
 wire \mod.pc[10] ;
 wire \mod.pc[11] ;
 wire \mod.pc[12] ;
 wire \mod.pc[13] ;
 wire \mod.pc[1] ;
 wire \mod.pc[2] ;
 wire \mod.pc[3] ;
 wire \mod.pc[4] ;
 wire \mod.pc[5] ;
 wire \mod.pc[6] ;
 wire \mod.pc[7] ;
 wire \mod.pc[8] ;
 wire \mod.pc[9] ;
 wire \mod.pc_1[0] ;
 wire \mod.pc_1[10] ;
 wire \mod.pc_1[11] ;
 wire \mod.pc_1[12] ;
 wire \mod.pc_1[13] ;
 wire \mod.pc_1[1] ;
 wire \mod.pc_1[2] ;
 wire \mod.pc_1[3] ;
 wire \mod.pc_1[4] ;
 wire \mod.pc_1[5] ;
 wire \mod.pc_1[6] ;
 wire \mod.pc_1[7] ;
 wire \mod.pc_1[8] ;
 wire \mod.pc_1[9] ;
 wire \mod.pc_2[0] ;
 wire \mod.pc_2[10] ;
 wire \mod.pc_2[11] ;
 wire \mod.pc_2[12] ;
 wire \mod.pc_2[13] ;
 wire \mod.pc_2[1] ;
 wire \mod.pc_2[2] ;
 wire \mod.pc_2[3] ;
 wire \mod.pc_2[4] ;
 wire \mod.pc_2[5] ;
 wire \mod.pc_2[6] ;
 wire \mod.pc_2[7] ;
 wire \mod.pc_2[8] ;
 wire \mod.pc_2[9] ;
 wire \mod.rd_3[0] ;
 wire \mod.rd_3[1] ;
 wire \mod.rd_3[2] ;
 wire \mod.rd_3[3] ;
 wire \mod.registers.r10[0] ;
 wire \mod.registers.r10[10] ;
 wire \mod.registers.r10[11] ;
 wire \mod.registers.r10[12] ;
 wire \mod.registers.r10[13] ;
 wire \mod.registers.r10[14] ;
 wire \mod.registers.r10[15] ;
 wire \mod.registers.r10[1] ;
 wire \mod.registers.r10[2] ;
 wire \mod.registers.r10[3] ;
 wire \mod.registers.r10[4] ;
 wire \mod.registers.r10[5] ;
 wire \mod.registers.r10[6] ;
 wire \mod.registers.r10[7] ;
 wire \mod.registers.r10[8] ;
 wire \mod.registers.r10[9] ;
 wire \mod.registers.r11[0] ;
 wire \mod.registers.r11[10] ;
 wire \mod.registers.r11[11] ;
 wire \mod.registers.r11[12] ;
 wire \mod.registers.r11[13] ;
 wire \mod.registers.r11[14] ;
 wire \mod.registers.r11[15] ;
 wire \mod.registers.r11[1] ;
 wire \mod.registers.r11[2] ;
 wire \mod.registers.r11[3] ;
 wire \mod.registers.r11[4] ;
 wire \mod.registers.r11[5] ;
 wire \mod.registers.r11[6] ;
 wire \mod.registers.r11[7] ;
 wire \mod.registers.r11[8] ;
 wire \mod.registers.r11[9] ;
 wire \mod.registers.r12[0] ;
 wire \mod.registers.r12[10] ;
 wire \mod.registers.r12[11] ;
 wire \mod.registers.r12[12] ;
 wire \mod.registers.r12[13] ;
 wire \mod.registers.r12[14] ;
 wire \mod.registers.r12[15] ;
 wire \mod.registers.r12[1] ;
 wire \mod.registers.r12[2] ;
 wire \mod.registers.r12[3] ;
 wire \mod.registers.r12[4] ;
 wire \mod.registers.r12[5] ;
 wire \mod.registers.r12[6] ;
 wire \mod.registers.r12[7] ;
 wire \mod.registers.r12[8] ;
 wire \mod.registers.r12[9] ;
 wire \mod.registers.r13[0] ;
 wire \mod.registers.r13[10] ;
 wire \mod.registers.r13[11] ;
 wire \mod.registers.r13[12] ;
 wire \mod.registers.r13[13] ;
 wire \mod.registers.r13[14] ;
 wire \mod.registers.r13[15] ;
 wire \mod.registers.r13[1] ;
 wire \mod.registers.r13[2] ;
 wire \mod.registers.r13[3] ;
 wire \mod.registers.r13[4] ;
 wire \mod.registers.r13[5] ;
 wire \mod.registers.r13[6] ;
 wire \mod.registers.r13[7] ;
 wire \mod.registers.r13[8] ;
 wire \mod.registers.r13[9] ;
 wire \mod.registers.r14[0] ;
 wire \mod.registers.r14[10] ;
 wire \mod.registers.r14[11] ;
 wire \mod.registers.r14[12] ;
 wire \mod.registers.r14[13] ;
 wire \mod.registers.r14[14] ;
 wire \mod.registers.r14[15] ;
 wire \mod.registers.r14[1] ;
 wire \mod.registers.r14[2] ;
 wire \mod.registers.r14[3] ;
 wire \mod.registers.r14[4] ;
 wire \mod.registers.r14[5] ;
 wire \mod.registers.r14[6] ;
 wire \mod.registers.r14[7] ;
 wire \mod.registers.r14[8] ;
 wire \mod.registers.r14[9] ;
 wire \mod.registers.r15[0] ;
 wire \mod.registers.r15[10] ;
 wire \mod.registers.r15[11] ;
 wire \mod.registers.r15[12] ;
 wire \mod.registers.r15[13] ;
 wire \mod.registers.r15[14] ;
 wire \mod.registers.r15[15] ;
 wire \mod.registers.r15[1] ;
 wire \mod.registers.r15[2] ;
 wire \mod.registers.r15[3] ;
 wire \mod.registers.r15[4] ;
 wire \mod.registers.r15[5] ;
 wire \mod.registers.r15[6] ;
 wire \mod.registers.r15[7] ;
 wire \mod.registers.r15[8] ;
 wire \mod.registers.r15[9] ;
 wire \mod.registers.r1[0] ;
 wire \mod.registers.r1[10] ;
 wire \mod.registers.r1[11] ;
 wire \mod.registers.r1[12] ;
 wire \mod.registers.r1[13] ;
 wire \mod.registers.r1[14] ;
 wire \mod.registers.r1[15] ;
 wire \mod.registers.r1[1] ;
 wire \mod.registers.r1[2] ;
 wire \mod.registers.r1[3] ;
 wire \mod.registers.r1[4] ;
 wire \mod.registers.r1[5] ;
 wire \mod.registers.r1[6] ;
 wire \mod.registers.r1[7] ;
 wire \mod.registers.r1[8] ;
 wire \mod.registers.r1[9] ;
 wire \mod.registers.r2[0] ;
 wire \mod.registers.r2[10] ;
 wire \mod.registers.r2[11] ;
 wire \mod.registers.r2[12] ;
 wire \mod.registers.r2[13] ;
 wire \mod.registers.r2[14] ;
 wire \mod.registers.r2[15] ;
 wire \mod.registers.r2[1] ;
 wire \mod.registers.r2[2] ;
 wire \mod.registers.r2[3] ;
 wire \mod.registers.r2[4] ;
 wire \mod.registers.r2[5] ;
 wire \mod.registers.r2[6] ;
 wire \mod.registers.r2[7] ;
 wire \mod.registers.r2[8] ;
 wire \mod.registers.r2[9] ;
 wire \mod.registers.r3[0] ;
 wire \mod.registers.r3[10] ;
 wire \mod.registers.r3[11] ;
 wire \mod.registers.r3[12] ;
 wire \mod.registers.r3[13] ;
 wire \mod.registers.r3[14] ;
 wire \mod.registers.r3[15] ;
 wire \mod.registers.r3[1] ;
 wire \mod.registers.r3[2] ;
 wire \mod.registers.r3[3] ;
 wire \mod.registers.r3[4] ;
 wire \mod.registers.r3[5] ;
 wire \mod.registers.r3[6] ;
 wire \mod.registers.r3[7] ;
 wire \mod.registers.r3[8] ;
 wire \mod.registers.r3[9] ;
 wire \mod.registers.r4[0] ;
 wire \mod.registers.r4[10] ;
 wire \mod.registers.r4[11] ;
 wire \mod.registers.r4[12] ;
 wire \mod.registers.r4[13] ;
 wire \mod.registers.r4[14] ;
 wire \mod.registers.r4[15] ;
 wire \mod.registers.r4[1] ;
 wire \mod.registers.r4[2] ;
 wire \mod.registers.r4[3] ;
 wire \mod.registers.r4[4] ;
 wire \mod.registers.r4[5] ;
 wire \mod.registers.r4[6] ;
 wire \mod.registers.r4[7] ;
 wire \mod.registers.r4[8] ;
 wire \mod.registers.r4[9] ;
 wire \mod.registers.r5[0] ;
 wire \mod.registers.r5[10] ;
 wire \mod.registers.r5[11] ;
 wire \mod.registers.r5[12] ;
 wire \mod.registers.r5[13] ;
 wire \mod.registers.r5[14] ;
 wire \mod.registers.r5[15] ;
 wire \mod.registers.r5[1] ;
 wire \mod.registers.r5[2] ;
 wire \mod.registers.r5[3] ;
 wire \mod.registers.r5[4] ;
 wire \mod.registers.r5[5] ;
 wire \mod.registers.r5[6] ;
 wire \mod.registers.r5[7] ;
 wire \mod.registers.r5[8] ;
 wire \mod.registers.r5[9] ;
 wire \mod.registers.r6[0] ;
 wire \mod.registers.r6[10] ;
 wire \mod.registers.r6[11] ;
 wire \mod.registers.r6[12] ;
 wire \mod.registers.r6[13] ;
 wire \mod.registers.r6[14] ;
 wire \mod.registers.r6[15] ;
 wire \mod.registers.r6[1] ;
 wire \mod.registers.r6[2] ;
 wire \mod.registers.r6[3] ;
 wire \mod.registers.r6[4] ;
 wire \mod.registers.r6[5] ;
 wire \mod.registers.r6[6] ;
 wire \mod.registers.r6[7] ;
 wire \mod.registers.r6[8] ;
 wire \mod.registers.r6[9] ;
 wire \mod.registers.r7[0] ;
 wire \mod.registers.r7[10] ;
 wire \mod.registers.r7[11] ;
 wire \mod.registers.r7[12] ;
 wire \mod.registers.r7[13] ;
 wire \mod.registers.r7[14] ;
 wire \mod.registers.r7[15] ;
 wire \mod.registers.r7[1] ;
 wire \mod.registers.r7[2] ;
 wire \mod.registers.r7[3] ;
 wire \mod.registers.r7[4] ;
 wire \mod.registers.r7[5] ;
 wire \mod.registers.r7[6] ;
 wire \mod.registers.r7[7] ;
 wire \mod.registers.r7[8] ;
 wire \mod.registers.r7[9] ;
 wire \mod.registers.r8[0] ;
 wire \mod.registers.r8[10] ;
 wire \mod.registers.r8[11] ;
 wire \mod.registers.r8[12] ;
 wire \mod.registers.r8[13] ;
 wire \mod.registers.r8[14] ;
 wire \mod.registers.r8[15] ;
 wire \mod.registers.r8[1] ;
 wire \mod.registers.r8[2] ;
 wire \mod.registers.r8[3] ;
 wire \mod.registers.r8[4] ;
 wire \mod.registers.r8[5] ;
 wire \mod.registers.r8[6] ;
 wire \mod.registers.r8[7] ;
 wire \mod.registers.r8[8] ;
 wire \mod.registers.r8[9] ;
 wire \mod.registers.r9[0] ;
 wire \mod.registers.r9[10] ;
 wire \mod.registers.r9[11] ;
 wire \mod.registers.r9[12] ;
 wire \mod.registers.r9[13] ;
 wire \mod.registers.r9[14] ;
 wire \mod.registers.r9[15] ;
 wire \mod.registers.r9[1] ;
 wire \mod.registers.r9[2] ;
 wire \mod.registers.r9[3] ;
 wire \mod.registers.r9[4] ;
 wire \mod.registers.r9[5] ;
 wire \mod.registers.r9[6] ;
 wire \mod.registers.r9[7] ;
 wire \mod.registers.r9[8] ;
 wire \mod.registers.r9[9] ;
 wire \mod.ri_3 ;
 wire \mod.valid0 ;
 wire \mod.valid1 ;
 wire \mod.valid2 ;
 wire \mod.valid_out3 ;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net347;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net348;
 wire net376;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3264_ (.I(\mod.des.des_counter[0] ),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3265_ (.I(\mod.des.des_counter[1] ),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3266_ (.A1(_0000_),
    .A2(_3120_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3267_ (.A1(net184),
    .A2(_3121_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(_3122_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3269_ (.A1(\mod.des.des_counter[0] ),
    .A2(_3120_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3270_ (.A1(_0000_),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3271_ (.A1(_3123_),
    .A2(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3272_ (.I(_3125_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3273_ (.I(_3126_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3274_ (.A1(\mod.des.des_counter[2] ),
    .A2(_3121_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3275_ (.I(_3127_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3276_ (.I(\mod.instr_2[17] ),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3277_ (.I(\mod.instr_2[16] ),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3278_ (.I(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3279_ (.I(\mod.instr_2[15] ),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3280_ (.I(\mod.instr_2[14] ),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3281_ (.A1(_3131_),
    .A2(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3282_ (.A1(_3128_),
    .A2(_3130_),
    .A3(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3283_ (.I(_3134_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3284_ (.I(\mod.instr_2[17] ),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3285_ (.A1(_3136_),
    .A2(\mod.instr_2[16] ),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3286_ (.A1(_3133_),
    .A2(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3287_ (.I(_3138_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3288_ (.A1(\mod.registers.r7[0] ),
    .A2(_3135_),
    .B1(_3139_),
    .B2(\mod.registers.r3[0] ),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3289_ (.I(_3136_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3290_ (.A1(_3131_),
    .A2(_3132_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3291_ (.A1(_3141_),
    .A2(_3130_),
    .A3(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3292_ (.I(_3143_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3293_ (.I(\mod.instr_2[15] ),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3294_ (.I(\mod.instr_2[14] ),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3295_ (.I(_3146_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3296_ (.A1(_3145_),
    .A2(_3147_),
    .A3(_3137_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(_3148_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3298_ (.A1(\mod.registers.r4[0] ),
    .A2(_3144_),
    .B1(_3149_),
    .B2(\mod.registers.r1[0] ),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3299_ (.A1(_3140_),
    .A2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3300_ (.I(\mod.instr_2[15] ),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3301_ (.I(_3132_),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3302_ (.A1(_3128_),
    .A2(_3130_),
    .A3(_3152_),
    .A4(_3153_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3303_ (.A1(_3128_),
    .A2(_3129_),
    .A3(_3131_),
    .A4(_3146_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3304_ (.A1(_3152_),
    .A2(_3153_),
    .A3(_3137_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3305_ (.A1(\mod.registers.r6[0] ),
    .A2(_3154_),
    .B1(_3155_),
    .B2(\mod.registers.r5[0] ),
    .C1(_3156_),
    .C2(\mod.registers.r2[0] ),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3306_ (.I(\mod.instr_2[17] ),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3307_ (.I(_3158_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3308_ (.I(\mod.instr_2[16] ),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3309_ (.A1(_3159_),
    .A2(_3160_),
    .A3(_3152_),
    .A4(_3153_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3310_ (.I(\mod.instr_2[16] ),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3311_ (.A1(_3158_),
    .A2(_3162_),
    .A3(_3145_),
    .A4(_3147_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3312_ (.A1(\mod.registers.r10[0] ),
    .A2(_3161_),
    .B1(_3163_),
    .B2(\mod.registers.r9[0] ),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3313_ (.A1(_3159_),
    .A2(_3160_),
    .A3(_3133_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3314_ (.I(_3165_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3315_ (.A1(_3159_),
    .A2(_3160_),
    .A3(_3142_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3316_ (.I(_3167_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3317_ (.A1(\mod.registers.r11[0] ),
    .A2(_3166_),
    .B1(_3168_),
    .B2(\mod.registers.r8[0] ),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(_3136_),
    .A2(_3162_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3319_ (.A1(_3145_),
    .A2(_3147_),
    .A3(_3170_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3320_ (.I(_3171_),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3321_ (.I(_3152_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3322_ (.I(_3132_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3323_ (.A1(_3173_),
    .A2(_3174_),
    .A3(_3170_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3324_ (.I(_3175_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3325_ (.I(\mod.registers.r12[0] ),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3326_ (.I(_3142_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3327_ (.I(_3170_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3328_ (.I(_3162_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3329_ (.I(_3131_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3330_ (.A1(_3141_),
    .A2(_3180_),
    .A3(_3181_),
    .A4(_3174_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3331_ (.I(\mod.registers.r15[0] ),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3332_ (.A1(_3177_),
    .A2(_3178_),
    .A3(_3179_),
    .B1(_3182_),
    .B2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3333_ (.A1(\mod.registers.r13[0] ),
    .A2(_3172_),
    .B1(_3176_),
    .B2(\mod.registers.r14[0] ),
    .C(_3184_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3334_ (.A1(_3157_),
    .A2(_3164_),
    .A3(_3169_),
    .A4(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3335_ (.I(_3123_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3336_ (.I(_3187_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3337_ (.A1(_3151_),
    .A2(_3186_),
    .B(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3338_ (.I(_3124_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3339_ (.I(\mod.funct3[2] ),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3340_ (.I(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3341_ (.I(\mod.funct3[1] ),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3342_ (.I(\mod.instr_2[2] ),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3343_ (.I(_3194_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3344_ (.I(\mod.instr_2[0] ),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3345_ (.I(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(_3195_),
    .A2(_3197_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3347_ (.I(\mod.instr_2[1] ),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3348_ (.I(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3349_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3350_ (.A1(_3200_),
    .A2(_3201_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3351_ (.I(_3202_),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3352_ (.I(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3353_ (.I(_3204_),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3354_ (.A1(_3193_),
    .A2(_3198_),
    .A3(_3205_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3355_ (.I(_3206_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3356_ (.A1(_3192_),
    .A2(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3357_ (.I(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3358_ (.I(_3209_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3359_ (.I(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3360_ (.I(_3193_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3361_ (.I(\mod.funct3[0] ),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3362_ (.A1(_3212_),
    .A2(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3363_ (.I(_3204_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3364_ (.A1(_3192_),
    .A2(_3214_),
    .B(_3215_),
    .C(_3198_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3365_ (.I(_3216_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3366_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3367_ (.A1(\mod.instr_2[1] ),
    .A2(_3218_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3368_ (.I(_3219_),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3369_ (.I(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3370_ (.I(_3221_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3371_ (.I(_3222_),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3372_ (.I(\mod.pc_2[0] ),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3373_ (.I(_3220_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3374_ (.I(_3225_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3375_ (.I(\mod.instr_2[13] ),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3376_ (.I(\mod.instr_2[12] ),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3377_ (.I(_3228_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3378_ (.I(\mod.instr_2[10] ),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3379_ (.A1(\mod.instr_2[11] ),
    .A2(_3230_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3380_ (.A1(_3227_),
    .A2(_3229_),
    .A3(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3381_ (.I(_3232_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3382_ (.I(_3233_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3383_ (.I(\mod.instr_2[11] ),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3384_ (.I(_3235_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3385_ (.I(_3230_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3386_ (.A1(_3227_),
    .A2(_3229_),
    .A3(_3236_),
    .A4(_3237_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3387_ (.I(_3238_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3388_ (.A1(\mod.registers.r8[0] ),
    .A2(_3234_),
    .B1(_3239_),
    .B2(\mod.registers.r10[0] ),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3389_ (.I(\mod.instr_2[13] ),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3390_ (.I(\mod.instr_2[12] ),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3391_ (.A1(_3241_),
    .A2(_3242_),
    .A3(_3236_),
    .A4(_3237_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3392_ (.I(_3243_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3393_ (.A1(\mod.instr_2[13] ),
    .A2(_3228_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3394_ (.A1(_3236_),
    .A2(_3237_),
    .A3(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3395_ (.I(_3246_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3396_ (.A1(\mod.registers.r6[0] ),
    .A2(_3244_),
    .B1(_3247_),
    .B2(\mod.registers.r14[0] ),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3397_ (.A1(_3241_),
    .A2(_3228_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3398_ (.A1(_3235_),
    .A2(_3230_),
    .A3(_3249_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3399_ (.I(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3400_ (.A1(\mod.instr_2[11] ),
    .A2(\mod.instr_2[10] ),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3401_ (.A1(_3227_),
    .A2(_3229_),
    .A3(_3252_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3402_ (.I(_3253_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3403_ (.I(_3254_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3404_ (.A1(\mod.registers.r2[0] ),
    .A2(_3251_),
    .B1(_3255_),
    .B2(\mod.registers.r11[0] ),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3405_ (.I(_3242_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3406_ (.A1(_3241_),
    .A2(_3257_),
    .A3(_3231_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3407_ (.I(_3258_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3408_ (.I(_3259_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3409_ (.I(_3219_),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3410_ (.I(_3261_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3411_ (.A1(\mod.registers.r4[0] ),
    .A2(_3260_),
    .B(_3262_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3412_ (.A1(_3240_),
    .A2(_3248_),
    .A3(_3256_),
    .A4(_3263_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3413_ (.I(\mod.instr_2[13] ),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3414_ (.I(\mod.instr_2[11] ),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3415_ (.I(\mod.instr_2[10] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3416_ (.A1(_0411_),
    .A2(_3242_),
    .A3(_0412_),
    .A4(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3417_ (.I(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3418_ (.A1(\mod.registers.r5[0] ),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3419_ (.A1(_0411_),
    .A2(_3257_),
    .A3(_3252_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3420_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(\mod.registers.r7[0] ),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3422_ (.I(_3227_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3423_ (.I(_3228_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3424_ (.A1(_0420_),
    .A2(_0421_),
    .A3(_0412_),
    .A4(_0413_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_3252_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3427_ (.A1(_3249_),
    .A2(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3429_ (.A1(\mod.registers.r9[0] ),
    .A2(_0423_),
    .B1(_0426_),
    .B2(\mod.registers.r3[0] ),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3430_ (.I(_0412_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3431_ (.I(_0413_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3432_ (.A1(_0428_),
    .A2(_0429_),
    .A3(_3249_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3433_ (.I(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3434_ (.A1(_0428_),
    .A2(_0429_),
    .A3(_3245_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3435_ (.I(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3436_ (.I(_3231_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3437_ (.I(_3245_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3438_ (.A1(_3241_),
    .A2(_3229_),
    .A3(_0412_),
    .A4(_3230_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3439_ (.A1(_3177_),
    .A2(_0434_),
    .A3(_0435_),
    .B1(_0436_),
    .B2(_3183_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3440_ (.A1(\mod.registers.r1[0] ),
    .A2(_0431_),
    .B1(_0433_),
    .B2(\mod.registers.r13[0] ),
    .C(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3441_ (.A1(_0416_),
    .A2(_0419_),
    .A3(_0427_),
    .A4(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3442_ (.A1(_3224_),
    .A2(_3226_),
    .B1(_0410_),
    .B2(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3443_ (.A1(_3199_),
    .A2(_3201_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3444_ (.I(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3445_ (.A1(_3200_),
    .A2(_3218_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3446_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3447_ (.I(_3174_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3448_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3449_ (.A1(\mod.funct3[2] ),
    .A2(_0446_),
    .B(_3201_),
    .C(\mod.instr_2[1] ),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3450_ (.I0(\mod.instr_2[3] ),
    .I1(_0445_),
    .S(_0447_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3451_ (.A1(_0444_),
    .A2(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3452_ (.A1(_0442_),
    .A2(_3151_),
    .A3(_3186_),
    .B(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3453_ (.I(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3454_ (.A1(_3223_),
    .A2(_0440_),
    .A3(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3455_ (.I(_3202_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3456_ (.A1(_3240_),
    .A2(_3248_),
    .A3(_3256_),
    .A4(_3263_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3457_ (.A1(_0416_),
    .A2(_0419_),
    .A3(_0427_),
    .A4(_0438_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3458_ (.A1(\mod.pc_2[0] ),
    .A2(_0453_),
    .B1(_0454_),
    .B2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3459_ (.I(_3225_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3460_ (.A1(_0457_),
    .A2(_0450_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3461_ (.I(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3462_ (.A1(_0456_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3463_ (.A1(_0452_),
    .A2(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3464_ (.I(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3465_ (.I(_3221_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3466_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3467_ (.A1(\mod.registers.r7[3] ),
    .A2(_3135_),
    .B1(_3138_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3468_ (.A1(\mod.registers.r4[3] ),
    .A2(_3143_),
    .B1(_3149_),
    .B2(\mod.registers.r1[3] ),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3469_ (.A1(_0465_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3470_ (.A1(\mod.registers.r6[3] ),
    .A2(_3154_),
    .B1(_3155_),
    .B2(\mod.registers.r5[3] ),
    .C1(_3156_),
    .C2(\mod.registers.r2[3] ),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3471_ (.A1(\mod.registers.r10[3] ),
    .A2(_3161_),
    .B1(_3163_),
    .B2(\mod.registers.r9[3] ),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3472_ (.A1(\mod.registers.r11[3] ),
    .A2(_3165_),
    .B1(_3167_),
    .B2(\mod.registers.r8[3] ),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3473_ (.I(\mod.registers.r12[3] ),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3474_ (.I(\mod.registers.r15[3] ),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3475_ (.A1(_0471_),
    .A2(_3178_),
    .A3(_3179_),
    .B1(_3182_),
    .B2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3476_ (.A1(\mod.registers.r13[3] ),
    .A2(_3172_),
    .B1(_3176_),
    .B2(\mod.registers.r14[3] ),
    .C(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3477_ (.A1(_0468_),
    .A2(_0469_),
    .A3(_0470_),
    .A4(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3478_ (.I(_3141_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3479_ (.I0(\mod.funct7[0] ),
    .I1(_0476_),
    .S(_0447_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3480_ (.A1(_0444_),
    .A2(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3481_ (.A1(_0442_),
    .A2(_0467_),
    .A3(_0475_),
    .B(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3482_ (.A1(_0464_),
    .A2(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3483_ (.I(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3484_ (.I(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3485_ (.I(_3250_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3486_ (.I(_0483_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3487_ (.I(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3488_ (.I(_3232_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3489_ (.I(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3490_ (.A1(\mod.registers.r2[15] ),
    .A2(_0485_),
    .B1(_0487_),
    .B2(\mod.registers.r8[15] ),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3491_ (.I(_0432_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3492_ (.I(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3493_ (.I(_3246_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3494_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3495_ (.A1(_0435_),
    .A2(_0424_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3496_ (.I(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3497_ (.I(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3498_ (.A1(\mod.registers.r13[15] ),
    .A2(_0490_),
    .B1(_0492_),
    .B2(\mod.registers.r14[15] ),
    .C1(\mod.registers.r15[15] ),
    .C2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3499_ (.I(_3255_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3500_ (.I(_3260_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3501_ (.A1(\mod.registers.r11[15] ),
    .A2(_0497_),
    .B1(_0498_),
    .B2(\mod.registers.r4[15] ),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3502_ (.A1(_0488_),
    .A2(_0496_),
    .A3(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3503_ (.I(_3244_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3504_ (.A1(_0434_),
    .A2(_0435_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3505_ (.I(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3506_ (.I(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3507_ (.A1(\mod.registers.r6[15] ),
    .A2(_0501_),
    .B1(_0504_),
    .B2(\mod.registers.r12[15] ),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3508_ (.I(_0422_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3509_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3510_ (.I(_3239_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3511_ (.A1(\mod.registers.r9[15] ),
    .A2(_0507_),
    .B1(_0508_),
    .B2(\mod.registers.r10[15] ),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3512_ (.I(_0430_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3513_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3514_ (.I(_0425_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3515_ (.I(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3516_ (.A1(\mod.registers.r1[15] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3517_ (.I(_0417_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3518_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3519_ (.I(_0414_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3520_ (.I(_0517_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3521_ (.A1(\mod.registers.r7[15] ),
    .A2(_0516_),
    .B1(_0518_),
    .B2(\mod.registers.r5[15] ),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3522_ (.A1(_0514_),
    .A2(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3523_ (.A1(_0500_),
    .A2(_0505_),
    .A3(_0509_),
    .A4(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3524_ (.A1(\mod.registers.r13[14] ),
    .A2(_0490_),
    .B1(_0498_),
    .B2(\mod.registers.r4[14] ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3525_ (.A1(\mod.registers.r6[14] ),
    .A2(_0501_),
    .B1(_0497_),
    .B2(\mod.registers.r11[14] ),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3526_ (.A1(\mod.registers.r1[14] ),
    .A2(_0511_),
    .B1(_0508_),
    .B2(\mod.registers.r10[14] ),
    .C1(\mod.registers.r14[14] ),
    .C2(_0492_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3527_ (.A1(_0522_),
    .A2(_0523_),
    .A3(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3528_ (.A1(\mod.registers.r9[14] ),
    .A2(_0507_),
    .B1(_0495_),
    .B2(\mod.registers.r15[14] ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3529_ (.A1(\mod.registers.r8[14] ),
    .A2(_0487_),
    .B1(_0504_),
    .B2(\mod.registers.r12[14] ),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3530_ (.A1(\mod.registers.r2[14] ),
    .A2(_0485_),
    .B1(_0513_),
    .B2(\mod.registers.r3[14] ),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3531_ (.A1(\mod.registers.r7[14] ),
    .A2(_0516_),
    .B1(_0518_),
    .B2(\mod.registers.r5[14] ),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3532_ (.A1(_0526_),
    .A2(_0527_),
    .A3(_0528_),
    .A4(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3533_ (.A1(_0525_),
    .A2(_0530_),
    .B(_3205_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3534_ (.A1(\mod.registers.r8[13] ),
    .A2(_0487_),
    .B1(_0508_),
    .B2(\mod.registers.r10[13] ),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3535_ (.A1(\mod.registers.r6[13] ),
    .A2(_0501_),
    .B1(_0492_),
    .B2(\mod.registers.r14[13] ),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3536_ (.A1(\mod.registers.r2[13] ),
    .A2(_0485_),
    .B1(_0497_),
    .B2(\mod.registers.r11[13] ),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3537_ (.I(_3262_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3538_ (.A1(\mod.registers.r4[13] ),
    .A2(_0498_),
    .B(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3539_ (.A1(_0532_),
    .A2(_0533_),
    .A3(_0534_),
    .A4(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3540_ (.A1(\mod.registers.r9[13] ),
    .A2(_0507_),
    .B1(_0513_),
    .B2(\mod.registers.r3[13] ),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3541_ (.A1(\mod.registers.r12[13] ),
    .A2(_0504_),
    .B1(_0495_),
    .B2(\mod.registers.r15[13] ),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3542_ (.A1(\mod.registers.r1[13] ),
    .A2(_0511_),
    .B1(_0490_),
    .B2(\mod.registers.r13[13] ),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3543_ (.A1(\mod.registers.r7[13] ),
    .A2(_0516_),
    .B1(_0518_),
    .B2(\mod.registers.r5[13] ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3544_ (.A1(_0538_),
    .A2(_0539_),
    .A3(_0540_),
    .A4(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3545_ (.A1(_0537_),
    .A2(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3546_ (.A1(\mod.pc_2[13] ),
    .A2(_3205_),
    .B(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3547_ (.A1(\mod.registers.r2[12] ),
    .A2(_0485_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3548_ (.A1(\mod.registers.r11[12] ),
    .A2(_0497_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3549_ (.A1(_0545_),
    .A2(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3550_ (.A1(\mod.registers.r8[12] ),
    .A2(_0487_),
    .B1(_0508_),
    .B2(\mod.registers.r10[12] ),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3551_ (.A1(\mod.registers.r6[12] ),
    .A2(_0501_),
    .B1(_0492_),
    .B2(\mod.registers.r14[12] ),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3552_ (.A1(_0548_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3553_ (.A1(\mod.registers.r4[12] ),
    .A2(_0498_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3554_ (.A1(_0453_),
    .A2(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3555_ (.A1(_0547_),
    .A2(_0550_),
    .A3(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3556_ (.A1(\mod.registers.r9[12] ),
    .A2(_0507_),
    .B1(_0513_),
    .B2(\mod.registers.r3[12] ),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3557_ (.A1(\mod.registers.r5[12] ),
    .A2(_0518_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3558_ (.A1(\mod.registers.r7[12] ),
    .A2(_0516_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3559_ (.A1(\mod.registers.r12[12] ),
    .A2(_0504_),
    .B1(_0495_),
    .B2(\mod.registers.r15[12] ),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3560_ (.A1(\mod.registers.r1[12] ),
    .A2(_0511_),
    .B1(_0490_),
    .B2(\mod.registers.r13[12] ),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3561_ (.A1(_0557_),
    .A2(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3562_ (.A1(_0554_),
    .A2(_0555_),
    .A3(_0556_),
    .A4(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3563_ (.A1(\mod.pc_2[12] ),
    .A2(_3215_),
    .B1(_0553_),
    .B2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3564_ (.A1(_3226_),
    .A2(_0450_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3565_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3566_ (.I(_0441_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3567_ (.I(_3143_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3568_ (.I(_3148_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3569_ (.A1(\mod.registers.r4[1] ),
    .A2(_0565_),
    .B1(_0566_),
    .B2(\mod.registers.r1[1] ),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3570_ (.I(_3155_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3571_ (.I(_3156_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3572_ (.A1(\mod.registers.r5[1] ),
    .A2(_0568_),
    .B1(_0569_),
    .B2(\mod.registers.r2[1] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3573_ (.A1(_0567_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3574_ (.I(_3154_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3575_ (.A1(\mod.registers.r7[1] ),
    .A2(_3135_),
    .B1(_0572_),
    .B2(\mod.registers.r6[1] ),
    .C1(_3139_),
    .C2(\mod.registers.r3[1] ),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3576_ (.I(_3167_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3577_ (.I(_3163_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3578_ (.A1(\mod.registers.r8[1] ),
    .A2(_0574_),
    .B1(_0575_),
    .B2(\mod.registers.r9[1] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3579_ (.I(_3165_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3580_ (.I(_3161_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3581_ (.A1(\mod.registers.r11[1] ),
    .A2(_0577_),
    .B1(_0578_),
    .B2(\mod.registers.r10[1] ),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(_3153_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3583_ (.A1(_3181_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3584_ (.A1(_3136_),
    .A2(_3162_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3585_ (.I(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3586_ (.A1(\mod.registers.r12[1] ),
    .A2(_0581_),
    .A3(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3587_ (.I(_3181_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3588_ (.I(_3147_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3589_ (.A1(_0585_),
    .A2(_0586_),
    .A3(\mod.registers.r14[1] ),
    .A4(_0582_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3590_ (.A1(_3173_),
    .A2(_0580_),
    .A3(\mod.registers.r13[1] ),
    .A4(_0582_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3591_ (.A1(_3128_),
    .A2(_3160_),
    .A3(_3145_),
    .A4(_3174_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3592_ (.A1(\mod.registers.r15[1] ),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3593_ (.A1(_0584_),
    .A2(_0587_),
    .A3(_0588_),
    .A4(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3594_ (.A1(_0573_),
    .A2(_0576_),
    .A3(_0579_),
    .A4(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3595_ (.A1(_0564_),
    .A2(_0571_),
    .A3(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3596_ (.I(_3202_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3597_ (.I(_0447_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3598_ (.I0(\mod.instr_2[4] ),
    .I1(_0585_),
    .S(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3599_ (.A1(_0444_),
    .A2(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3600_ (.A1(_0594_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_0593_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3602_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3603_ (.I0(_0521_),
    .I1(_0531_),
    .I2(_0544_),
    .I3(_0561_),
    .S0(_0563_),
    .S1(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3604_ (.I(_3238_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3605_ (.A1(\mod.registers.r8[11] ),
    .A2(_3234_),
    .B1(_0602_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3606_ (.I(_3243_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3607_ (.I(_3246_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3608_ (.A1(\mod.registers.r6[11] ),
    .A2(_0604_),
    .B1(_0605_),
    .B2(\mod.registers.r14[11] ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3609_ (.I(_0421_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3610_ (.I(_0428_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3611_ (.I(_3237_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3612_ (.A1(_0608_),
    .A2(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3613_ (.A1(_0420_),
    .A2(_0607_),
    .A3(\mod.registers.r4[11] ),
    .A4(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3614_ (.I(_0411_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3615_ (.A1(_0612_),
    .A2(_0421_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3616_ (.A1(_0608_),
    .A2(_0429_),
    .A3(\mod.registers.r2[11] ),
    .A4(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3617_ (.I(_0411_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_3257_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3619_ (.A1(_0428_),
    .A2(_0609_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3620_ (.A1(_0615_),
    .A2(_0616_),
    .A3(\mod.registers.r11[11] ),
    .A4(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3621_ (.A1(_3203_),
    .A2(_0611_),
    .A3(_0614_),
    .A4(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3622_ (.A1(_0603_),
    .A2(_0606_),
    .A3(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3623_ (.I(_0494_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3624_ (.A1(\mod.registers.r12[11] ),
    .A2(_0503_),
    .B1(_0621_),
    .B2(\mod.registers.r15[11] ),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3625_ (.I(_0422_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3626_ (.I(_0425_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3627_ (.A1(\mod.registers.r9[11] ),
    .A2(_0623_),
    .B1(_0624_),
    .B2(\mod.registers.r3[11] ),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3628_ (.A1(\mod.registers.r7[11] ),
    .A2(_0418_),
    .B1(_0415_),
    .B2(\mod.registers.r5[11] ),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3629_ (.I(_0432_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3630_ (.A1(\mod.registers.r1[11] ),
    .A2(_0510_),
    .B1(_0627_),
    .B2(\mod.registers.r13[11] ),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3631_ (.A1(_0622_),
    .A2(_0625_),
    .A3(_0626_),
    .A4(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3632_ (.A1(\mod.pc_2[11] ),
    .A2(_0453_),
    .B1(_0620_),
    .B2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3633_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3634_ (.I(_3238_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3635_ (.A1(\mod.registers.r8[10] ),
    .A2(_0486_),
    .B1(_0632_),
    .B2(\mod.registers.r10[10] ),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3636_ (.I(_3243_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3637_ (.A1(\mod.registers.r6[10] ),
    .A2(_0634_),
    .B1(_3247_),
    .B2(\mod.registers.r14[10] ),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3638_ (.I(_3254_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3639_ (.A1(\mod.registers.r2[10] ),
    .A2(_3251_),
    .B1(_0636_),
    .B2(\mod.registers.r11[10] ),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3640_ (.I(_3258_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3641_ (.I(_3261_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3642_ (.A1(\mod.registers.r4[10] ),
    .A2(_0638_),
    .B(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3643_ (.A1(_0633_),
    .A2(_0635_),
    .A3(_0637_),
    .A4(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3644_ (.A1(\mod.registers.r9[10] ),
    .A2(_0423_),
    .B1(_0426_),
    .B2(\mod.registers.r3[10] ),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3645_ (.I(_0502_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3646_ (.I(_0493_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3647_ (.A1(\mod.registers.r12[10] ),
    .A2(_0643_),
    .B1(_0644_),
    .B2(\mod.registers.r15[10] ),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3648_ (.A1(\mod.registers.r1[10] ),
    .A2(_0431_),
    .B1(_0433_),
    .B2(\mod.registers.r13[10] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3649_ (.A1(\mod.registers.r7[10] ),
    .A2(_0515_),
    .B1(_0517_),
    .B2(\mod.registers.r5[10] ),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3650_ (.A1(_0642_),
    .A2(_0645_),
    .A3(_0646_),
    .A4(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3651_ (.A1(\mod.pc_2[10] ),
    .A2(_3203_),
    .B1(_0641_),
    .B2(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3653_ (.A1(\mod.registers.r6[9] ),
    .A2(_0604_),
    .B1(_0605_),
    .B2(\mod.registers.r14[9] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3654_ (.A1(\mod.registers.r8[9] ),
    .A2(_3234_),
    .B1(_0602_),
    .B2(\mod.registers.r10[9] ),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3655_ (.A1(\mod.registers.r2[9] ),
    .A2(_0484_),
    .B1(_3255_),
    .B2(\mod.registers.r11[9] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3656_ (.A1(\mod.registers.r4[9] ),
    .A2(_3260_),
    .B(_3221_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3657_ (.A1(_0651_),
    .A2(_0652_),
    .A3(_0653_),
    .A4(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3658_ (.A1(\mod.registers.r7[9] ),
    .A2(_0418_),
    .B1(_0415_),
    .B2(\mod.registers.r5[9] ),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3659_ (.A1(\mod.registers.r9[9] ),
    .A2(_0623_),
    .B1(_0624_),
    .B2(\mod.registers.r3[9] ),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3660_ (.A1(\mod.registers.r12[9] ),
    .A2(_0503_),
    .B1(_0621_),
    .B2(\mod.registers.r15[9] ),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3661_ (.A1(\mod.registers.r1[9] ),
    .A2(_0510_),
    .B1(_0627_),
    .B2(\mod.registers.r13[9] ),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3662_ (.A1(_0656_),
    .A2(_0657_),
    .A3(_0658_),
    .A4(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3663_ (.A1(\mod.pc_2[9] ),
    .A2(_3204_),
    .B1(_0655_),
    .B2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3664_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3665_ (.I(\mod.pc_2[8] ),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3666_ (.A1(\mod.registers.r4[8] ),
    .A2(_3260_),
    .B1(_0621_),
    .B2(\mod.registers.r15[8] ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3667_ (.A1(\mod.registers.r6[8] ),
    .A2(_0604_),
    .B1(_0418_),
    .B2(\mod.registers.r7[8] ),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3668_ (.A1(_0612_),
    .A2(_3257_),
    .A3(\mod.registers.r11[8] ),
    .A4(_0617_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3669_ (.A1(_0612_),
    .A2(_0421_),
    .A3(\mod.registers.r12[8] ),
    .A4(_0610_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3670_ (.A1(_0612_),
    .A2(_0616_),
    .A3(\mod.registers.r8[8] ),
    .A4(_0610_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3671_ (.A1(_3202_),
    .A2(_0666_),
    .A3(_0667_),
    .A4(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3672_ (.A1(_0664_),
    .A2(_0665_),
    .A3(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3673_ (.A1(\mod.registers.r1[8] ),
    .A2(_0510_),
    .B1(_0624_),
    .B2(\mod.registers.r3[8] ),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3674_ (.A1(\mod.registers.r10[8] ),
    .A2(_0602_),
    .B1(_0627_),
    .B2(\mod.registers.r13[8] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3675_ (.A1(\mod.registers.r9[8] ),
    .A2(_0623_),
    .B1(_0605_),
    .B2(\mod.registers.r14[8] ),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3676_ (.A1(\mod.registers.r2[8] ),
    .A2(_0484_),
    .B1(_0415_),
    .B2(\mod.registers.r5[8] ),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3677_ (.A1(_0671_),
    .A2(_0672_),
    .A3(_0673_),
    .A4(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3678_ (.A1(_0663_),
    .A2(_3215_),
    .B1(_0670_),
    .B2(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3679_ (.I0(_0631_),
    .I1(_0650_),
    .I2(_0662_),
    .I3(_0676_),
    .S0(_0563_),
    .S1(_0600_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3680_ (.I(_0535_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3681_ (.I(_3134_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(_3138_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3683_ (.A1(\mod.registers.r7[2] ),
    .A2(_0679_),
    .B1(_0680_),
    .B2(\mod.registers.r3[2] ),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3684_ (.A1(\mod.registers.r4[2] ),
    .A2(_0565_),
    .B1(_0566_),
    .B2(\mod.registers.r1[2] ),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3685_ (.A1(_0681_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3686_ (.I(_3154_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3687_ (.A1(\mod.registers.r6[2] ),
    .A2(_0684_),
    .B1(_0568_),
    .B2(\mod.registers.r5[2] ),
    .C1(_0569_),
    .C2(\mod.registers.r2[2] ),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3688_ (.I(_3161_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3689_ (.A1(\mod.registers.r10[2] ),
    .A2(_0686_),
    .B1(_0575_),
    .B2(\mod.registers.r9[2] ),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3690_ (.A1(\mod.registers.r11[2] ),
    .A2(_0577_),
    .B1(_0574_),
    .B2(\mod.registers.r8[2] ),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3691_ (.I(_3171_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3692_ (.I(_3175_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3693_ (.I(\mod.registers.r12[2] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3694_ (.I(\mod.registers.r15[2] ),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3695_ (.A1(_0691_),
    .A2(_3178_),
    .A3(_3179_),
    .B1(_3182_),
    .B2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3696_ (.A1(\mod.registers.r13[2] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\mod.registers.r14[2] ),
    .C(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3697_ (.A1(_0685_),
    .A2(_0687_),
    .A3(_0688_),
    .A4(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3698_ (.I(_0443_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3699_ (.I(_3180_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3700_ (.I0(\mod.instr_2[5] ),
    .I1(_0697_),
    .S(_0595_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3701_ (.A1(_0696_),
    .A2(_0698_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3702_ (.A1(_0564_),
    .A2(_0683_),
    .A3(_0695_),
    .B(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3703_ (.A1(_0678_),
    .A2(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3704_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3705_ (.I0(_0601_),
    .I1(_0677_),
    .S(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3706_ (.A1(_0482_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3707_ (.I(_3226_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3708_ (.I(_0441_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3709_ (.A1(\mod.registers.r7[4] ),
    .A2(_0679_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3710_ (.A1(\mod.registers.r3[4] ),
    .A2(_0680_),
    .B1(_0566_),
    .B2(\mod.registers.r1[4] ),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3711_ (.A1(\mod.registers.r5[4] ),
    .A2(_0568_),
    .B1(_0574_),
    .B2(\mod.registers.r8[4] ),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3712_ (.I(_0589_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3713_ (.I(_3163_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3714_ (.A1(\mod.registers.r15[4] ),
    .A2(_0710_),
    .B1(_0711_),
    .B2(\mod.registers.r9[4] ),
    .C1(\mod.registers.r6[4] ),
    .C2(_0684_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3715_ (.A1(_0707_),
    .A2(_0708_),
    .A3(_0709_),
    .A4(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3716_ (.A1(\mod.registers.r2[4] ),
    .A2(_0569_),
    .B1(_3144_),
    .B2(\mod.registers.r4[4] ),
    .C1(\mod.registers.r10[4] ),
    .C2(_0686_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3717_ (.A1(_3142_),
    .A2(_3170_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3718_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3719_ (.A1(\mod.registers.r12[4] ),
    .A2(_0716_),
    .B1(_0690_),
    .B2(\mod.registers.r14[4] ),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3720_ (.A1(\mod.registers.r13[4] ),
    .A2(_0689_),
    .B1(_0577_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3721_ (.A1(_0714_),
    .A2(_0717_),
    .A3(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3722_ (.I0(\mod.funct7[1] ),
    .I1(\mod.funct7[0] ),
    .S(_0595_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3723_ (.A1(_0444_),
    .A2(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3724_ (.A1(_0706_),
    .A2(_0713_),
    .A3(_0719_),
    .B(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3725_ (.A1(_0705_),
    .A2(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3726_ (.A1(_0500_),
    .A2(_0505_),
    .A3(_0509_),
    .A4(_0520_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3727_ (.I(_3199_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3728_ (.I(_0446_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_0725_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3730_ (.I(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3731_ (.A1(_3191_),
    .A2(_0725_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3732_ (.A1(\mod.funct7[1] ),
    .A2(_3196_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3733_ (.A1(_3194_),
    .A2(_0729_),
    .A3(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3734_ (.A1(_0728_),
    .A2(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3735_ (.A1(_0724_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3736_ (.A1(_0723_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3737_ (.A1(_0705_),
    .A2(_0479_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3738_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3739_ (.I(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3740_ (.A1(_0464_),
    .A2(_0700_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3741_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3742_ (.I(\mod.pc_2[7] ),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3743_ (.A1(\mod.registers.r8[7] ),
    .A2(_3233_),
    .B1(_0632_),
    .B2(\mod.registers.r10[7] ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3744_ (.A1(\mod.registers.r6[7] ),
    .A2(_0634_),
    .B1(_0491_),
    .B2(\mod.registers.r14[7] ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3745_ (.A1(\mod.registers.r2[7] ),
    .A2(_0483_),
    .B1(_3254_),
    .B2(\mod.registers.r11[7] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3746_ (.A1(\mod.registers.r4[7] ),
    .A2(_3259_),
    .B(_3261_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3747_ (.A1(_0741_),
    .A2(_0742_),
    .A3(_0743_),
    .A4(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3748_ (.A1(\mod.registers.r12[7] ),
    .A2(_0502_),
    .B1(_0494_),
    .B2(\mod.registers.r15[7] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3749_ (.I(_0430_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3750_ (.A1(\mod.registers.r1[7] ),
    .A2(_0747_),
    .B1(_0489_),
    .B2(\mod.registers.r13[7] ),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3751_ (.A1(\mod.registers.r9[7] ),
    .A2(_0506_),
    .B1(_0512_),
    .B2(\mod.registers.r3[7] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3752_ (.I(_0417_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3753_ (.I(_0414_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3754_ (.A1(\mod.registers.r7[7] ),
    .A2(_0750_),
    .B1(_0751_),
    .B2(\mod.registers.r5[7] ),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3755_ (.A1(_0746_),
    .A2(_0748_),
    .A3(_0749_),
    .A4(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3756_ (.A1(_0745_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3757_ (.A1(_0740_),
    .A2(_3225_),
    .B(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3758_ (.A1(\mod.registers.r8[6] ),
    .A2(_3234_),
    .B1(_0602_),
    .B2(\mod.registers.r10[6] ),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3759_ (.A1(\mod.registers.r6[6] ),
    .A2(_0604_),
    .B1(_0605_),
    .B2(\mod.registers.r14[6] ),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3760_ (.A1(\mod.registers.r2[6] ),
    .A2(_0484_),
    .B1(_3255_),
    .B2(\mod.registers.r11[6] ),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3761_ (.A1(\mod.registers.r4[6] ),
    .A2(_0638_),
    .B(_3262_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3762_ (.A1(_0756_),
    .A2(_0757_),
    .A3(_0758_),
    .A4(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3763_ (.A1(\mod.registers.r12[6] ),
    .A2(_0503_),
    .B1(_0621_),
    .B2(\mod.registers.r15[6] ),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3764_ (.A1(\mod.registers.r1[6] ),
    .A2(_0431_),
    .B1(_0627_),
    .B2(\mod.registers.r13[6] ),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3765_ (.A1(\mod.registers.r9[6] ),
    .A2(_0623_),
    .B1(_0624_),
    .B2(\mod.registers.r3[6] ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3766_ (.A1(\mod.registers.r7[6] ),
    .A2(_0515_),
    .B1(_0517_),
    .B2(\mod.registers.r5[6] ),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3767_ (.A1(_0761_),
    .A2(_0762_),
    .A3(_0763_),
    .A4(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3768_ (.A1(\mod.pc_2[6] ),
    .A2(_0594_),
    .B1(_0760_),
    .B2(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3769_ (.I(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(\mod.pc_2[5] ),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3771_ (.I(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3772_ (.A1(\mod.registers.r8[5] ),
    .A2(_3233_),
    .B1(_0632_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3773_ (.A1(\mod.registers.r6[5] ),
    .A2(_0634_),
    .B1(_0491_),
    .B2(\mod.registers.r14[5] ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3774_ (.A1(\mod.registers.r2[5] ),
    .A2(_0483_),
    .B1(_3254_),
    .B2(\mod.registers.r11[5] ),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3775_ (.A1(\mod.registers.r4[5] ),
    .A2(_3259_),
    .B(_3220_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3776_ (.A1(_0770_),
    .A2(_0771_),
    .A3(_0772_),
    .A4(_0773_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3777_ (.A1(\mod.registers.r9[5] ),
    .A2(_0506_),
    .B1(_0512_),
    .B2(\mod.registers.r3[5] ),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3778_ (.A1(\mod.registers.r12[5] ),
    .A2(_0502_),
    .B1(_0494_),
    .B2(\mod.registers.r15[5] ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3779_ (.A1(\mod.registers.r7[5] ),
    .A2(_0750_),
    .B1(_0751_),
    .B2(\mod.registers.r5[5] ),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3780_ (.A1(\mod.registers.r1[5] ),
    .A2(_0747_),
    .B1(_0489_),
    .B2(\mod.registers.r13[5] ),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3781_ (.A1(_0775_),
    .A2(_0776_),
    .A3(_0777_),
    .A4(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3782_ (.A1(_0769_),
    .A2(_0678_),
    .B1(_0774_),
    .B2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3783_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3784_ (.A1(\mod.registers.r5[4] ),
    .A2(_0751_),
    .B1(_0644_),
    .B2(\mod.registers.r15[4] ),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3785_ (.A1(\mod.registers.r9[4] ),
    .A2(_0506_),
    .B1(_0636_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3786_ (.A1(\mod.registers.r2[4] ),
    .A2(_3251_),
    .B(_0639_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3787_ (.A1(\mod.registers.r12[4] ),
    .A2(_0643_),
    .B1(_3247_),
    .B2(\mod.registers.r14[4] ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3788_ (.A1(_0782_),
    .A2(_0783_),
    .A3(_0784_),
    .A4(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3789_ (.A1(\mod.registers.r10[4] ),
    .A2(_3239_),
    .B1(_0638_),
    .B2(\mod.registers.r4[4] ),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3790_ (.A1(\mod.registers.r8[4] ),
    .A2(_0486_),
    .B1(_0747_),
    .B2(\mod.registers.r1[4] ),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3791_ (.A1(\mod.registers.r13[4] ),
    .A2(_0433_),
    .B1(_0512_),
    .B2(\mod.registers.r3[4] ),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3792_ (.A1(\mod.registers.r6[4] ),
    .A2(_3244_),
    .B1(_0750_),
    .B2(\mod.registers.r7[4] ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3793_ (.A1(_0787_),
    .A2(_0788_),
    .A3(_0789_),
    .A4(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3794_ (.A1(_0786_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3795_ (.A1(\mod.pc_2[4] ),
    .A2(_3204_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3796_ (.A1(_0792_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3797_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3798_ (.I(_0562_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3799_ (.I(_0599_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3800_ (.I0(_0755_),
    .I1(_0767_),
    .I2(_0781_),
    .I3(_0795_),
    .S0(_0796_),
    .S1(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3801_ (.I(\mod.pc_2[3] ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3802_ (.A1(\mod.registers.r8[3] ),
    .A2(_3232_),
    .B1(_3238_),
    .B2(\mod.registers.r10[3] ),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3803_ (.A1(\mod.registers.r6[3] ),
    .A2(_3243_),
    .B1(_3246_),
    .B2(\mod.registers.r14[3] ),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3804_ (.A1(\mod.registers.r2[3] ),
    .A2(_3250_),
    .B1(_3253_),
    .B2(\mod.registers.r11[3] ),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3805_ (.A1(\mod.registers.r4[3] ),
    .A2(_3258_),
    .B(_3261_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3806_ (.A1(_0800_),
    .A2(_0801_),
    .A3(_0802_),
    .A4(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3807_ (.A1(\mod.registers.r5[3] ),
    .A2(_0414_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(\mod.registers.r7[3] ),
    .A2(_0417_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3809_ (.A1(\mod.registers.r9[3] ),
    .A2(_0422_),
    .B1(_0425_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3810_ (.A1(_0471_),
    .A2(_3231_),
    .A3(_0435_),
    .B1(_0436_),
    .B2(_0472_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3811_ (.A1(\mod.registers.r1[3] ),
    .A2(_0430_),
    .B1(_0432_),
    .B2(\mod.registers.r13[3] ),
    .C(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3812_ (.A1(_0805_),
    .A2(_0806_),
    .A3(_0807_),
    .A4(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3813_ (.A1(_0799_),
    .A2(_3262_),
    .B1(_0804_),
    .B2(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3814_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3815_ (.I(\mod.pc_2[2] ),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3816_ (.A1(\mod.registers.r8[2] ),
    .A2(_3233_),
    .B1(_0632_),
    .B2(\mod.registers.r10[2] ),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3817_ (.A1(\mod.registers.r6[2] ),
    .A2(_0634_),
    .B1(_0491_),
    .B2(\mod.registers.r14[2] ),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3818_ (.A1(\mod.registers.r2[2] ),
    .A2(_0483_),
    .B1(_0636_),
    .B2(\mod.registers.r11[2] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3819_ (.A1(\mod.registers.r4[2] ),
    .A2(_3259_),
    .B(_0639_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3820_ (.A1(_0814_),
    .A2(_0815_),
    .A3(_0816_),
    .A4(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3821_ (.A1(\mod.registers.r9[2] ),
    .A2(_0423_),
    .B1(_0426_),
    .B2(\mod.registers.r3[2] ),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3822_ (.A1(\mod.registers.r12[2] ),
    .A2(_0643_),
    .B1(_0644_),
    .B2(\mod.registers.r15[2] ),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3823_ (.A1(\mod.registers.r7[2] ),
    .A2(_0750_),
    .B1(_0751_),
    .B2(\mod.registers.r5[2] ),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3824_ (.A1(\mod.registers.r1[2] ),
    .A2(_0747_),
    .B1(_0489_),
    .B2(\mod.registers.r13[2] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3825_ (.A1(_0819_),
    .A2(_0820_),
    .A3(_0821_),
    .A4(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3826_ (.A1(_0813_),
    .A2(_3222_),
    .B1(_0818_),
    .B2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3827_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3828_ (.I(_0562_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3829_ (.I0(_0812_),
    .I1(_0825_),
    .S(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3830_ (.I(_0738_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3831_ (.A1(_0600_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3832_ (.I(\mod.pc_2[1] ),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3833_ (.A1(\mod.registers.r8[1] ),
    .A2(_0486_),
    .B1(_0433_),
    .B2(\mod.registers.r13[1] ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3834_ (.A1(\mod.registers.r6[1] ),
    .A2(_3244_),
    .B1(_0643_),
    .B2(\mod.registers.r12[1] ),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3835_ (.A1(\mod.registers.r2[1] ),
    .A2(_3251_),
    .B1(_0431_),
    .B2(\mod.registers.r1[1] ),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3836_ (.A1(\mod.registers.r4[1] ),
    .A2(_0638_),
    .B(_0639_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3837_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0833_),
    .A4(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3838_ (.A1(\mod.registers.r3[1] ),
    .A2(_0426_),
    .B1(_0644_),
    .B2(\mod.registers.r15[1] ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3839_ (.A1(\mod.registers.r11[1] ),
    .A2(_0636_),
    .B1(_3247_),
    .B2(\mod.registers.r14[1] ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3840_ (.A1(\mod.registers.r7[1] ),
    .A2(_0515_),
    .B1(_0517_),
    .B2(\mod.registers.r5[1] ),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3841_ (.A1(\mod.registers.r9[1] ),
    .A2(_0423_),
    .B1(_3239_),
    .B2(\mod.registers.r10[1] ),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3842_ (.A1(_0836_),
    .A2(_0837_),
    .A3(_0838_),
    .A4(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3843_ (.A1(_0830_),
    .A2(_0463_),
    .B1(_0835_),
    .B2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3844_ (.I(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3845_ (.I0(_0842_),
    .I1(_0440_),
    .S(_0826_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3846_ (.A1(_0706_),
    .A2(_0571_),
    .A3(_0592_),
    .B(_0597_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3847_ (.A1(_0463_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3848_ (.I(_0845_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3849_ (.A1(_0846_),
    .A2(_0828_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3850_ (.A1(_0739_),
    .A2(_0798_),
    .B1(_0827_),
    .B2(_0829_),
    .C1(_0843_),
    .C2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3851_ (.A1(_0737_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3852_ (.I(_3191_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3853_ (.I(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3854_ (.I(\mod.funct3[0] ),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3855_ (.I(_0678_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3856_ (.A1(_3193_),
    .A2(_0726_),
    .A3(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3857_ (.A1(_0852_),
    .A2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3858_ (.A1(_0851_),
    .A2(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3859_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3860_ (.A1(_0704_),
    .A2(_0734_),
    .A3(_0849_),
    .B(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3861_ (.A1(_0850_),
    .A2(_3213_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3862_ (.A1(_3206_),
    .A2(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3863_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3864_ (.I(_0563_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3865_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3866_ (.A1(_0456_),
    .A2(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3867_ (.A1(_0850_),
    .A2(_0852_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3868_ (.A1(_0865_),
    .A2(_3206_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3869_ (.A1(_0457_),
    .A2(_0456_),
    .A3(_0451_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3870_ (.A1(_0866_),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3871_ (.I(_3216_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3872_ (.A1(_0861_),
    .A2(_0864_),
    .B(_0868_),
    .C(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3873_ (.A1(_0851_),
    .A2(_0852_),
    .A3(_0854_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3874_ (.A1(_0736_),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3875_ (.A1(_0847_),
    .A2(_0460_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3876_ (.I(_3213_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3877_ (.A1(_0850_),
    .A2(_0874_),
    .A3(_0854_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3878_ (.A1(_3208_),
    .A2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3879_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0461_),
    .B2(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3880_ (.A1(_0870_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3881_ (.A1(_3217_),
    .A2(_0462_),
    .B1(_0858_),
    .B2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_3211_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3883_ (.I(_0853_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3884_ (.I(_0521_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3885_ (.A1(_0881_),
    .A2(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3886_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3887_ (.I(_3159_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3888_ (.A1(_0726_),
    .A2(_0441_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3889_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3890_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3891_ (.I(\mod.funct7[2] ),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3892_ (.A1(_0889_),
    .A2(_0887_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3893_ (.A1(_0885_),
    .A2(_0888_),
    .B(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3894_ (.I(_3135_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3895_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3896_ (.I(_0578_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3897_ (.I(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3898_ (.I(_3155_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3899_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3900_ (.I(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3901_ (.I(_3139_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3902_ (.I(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3903_ (.A1(\mod.registers.r5[15] ),
    .A2(_0898_),
    .B1(_0900_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3904_ (.I(_0572_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3905_ (.I(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3906_ (.I(_0715_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3907_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3908_ (.A1(\mod.registers.r6[15] ),
    .A2(_0903_),
    .B1(_0905_),
    .B2(\mod.registers.r12[15] ),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3909_ (.I(_3144_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3910_ (.I(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3911_ (.I(_3168_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3912_ (.I(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3913_ (.A1(\mod.registers.r4[15] ),
    .A2(_0908_),
    .B1(_0910_),
    .B2(\mod.registers.r8[15] ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3914_ (.A1(_0901_),
    .A2(_0906_),
    .A3(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3915_ (.A1(\mod.registers.r7[15] ),
    .A2(_0893_),
    .B1(_0895_),
    .B2(\mod.registers.r10[15] ),
    .C(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3916_ (.I(_0696_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3917_ (.I(_3165_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3918_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3919_ (.I(_3176_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3920_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3921_ (.I(_0589_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3922_ (.I(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3923_ (.A1(\mod.registers.r11[15] ),
    .A2(_0916_),
    .B1(_0918_),
    .B2(\mod.registers.r14[15] ),
    .C1(\mod.registers.r15[15] ),
    .C2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3924_ (.I(_3156_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3925_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3926_ (.I(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3927_ (.I(_3149_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3928_ (.I(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3929_ (.A1(\mod.registers.r2[15] ),
    .A2(_0924_),
    .B1(_0926_),
    .B2(\mod.registers.r1[15] ),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_3172_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3932_ (.I(_0711_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3933_ (.I(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3934_ (.A1(\mod.registers.r13[15] ),
    .A2(_0929_),
    .B1(_0931_),
    .B2(\mod.registers.r9[15] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3935_ (.A1(_0914_),
    .A2(_0921_),
    .A3(_0927_),
    .A4(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3936_ (.I(_3218_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3937_ (.A1(_0889_),
    .A2(_0934_),
    .B(_0725_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3938_ (.A1(_0913_),
    .A2(_0933_),
    .B(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3939_ (.A1(_0881_),
    .A2(_0891_),
    .B(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_0724_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3941_ (.A1(_3215_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3942_ (.A1(_0939_),
    .A2(_0937_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(_0938_),
    .A2(_0936_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3944_ (.A1(_0940_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3945_ (.I(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3946_ (.I(_0726_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3947_ (.I(_3192_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3948_ (.A1(_0945_),
    .A2(_3214_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3949_ (.A1(_0944_),
    .A2(_0881_),
    .A3(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3951_ (.A1(\mod.registers.r5[7] ),
    .A2(_0896_),
    .B1(_0578_),
    .B2(\mod.registers.r10[7] ),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3952_ (.A1(\mod.registers.r15[7] ),
    .A2(_0589_),
    .B1(_0711_),
    .B2(\mod.registers.r9[7] ),
    .C1(\mod.registers.r6[7] ),
    .C2(_0572_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3953_ (.A1(\mod.registers.r2[7] ),
    .A2(_0922_),
    .B1(_3166_),
    .B2(\mod.registers.r11[7] ),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3954_ (.A1(_0949_),
    .A2(_0950_),
    .A3(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3955_ (.A1(\mod.registers.r12[7] ),
    .A2(_0716_),
    .B1(_0689_),
    .B2(\mod.registers.r13[7] ),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3956_ (.A1(\mod.registers.r1[7] ),
    .A2(_3149_),
    .B1(_3168_),
    .B2(\mod.registers.r8[7] ),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3957_ (.A1(\mod.registers.r3[7] ),
    .A2(_0680_),
    .B1(_3144_),
    .B2(\mod.registers.r4[7] ),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3958_ (.A1(\mod.registers.r7[7] ),
    .A2(_0679_),
    .B1(_0690_),
    .B2(\mod.registers.r14[7] ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3959_ (.A1(_0953_),
    .A2(_0954_),
    .A3(_0955_),
    .A4(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3960_ (.A1(\mod.funct7[2] ),
    .A2(_0443_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3961_ (.A1(_3220_),
    .A2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3962_ (.A1(_0442_),
    .A2(_0952_),
    .A3(_0957_),
    .B(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3963_ (.I0(_0698_),
    .I1(_3191_),
    .S(_0886_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3964_ (.A1(_3225_),
    .A2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3965_ (.A1(_0960_),
    .A2(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3966_ (.A1(_0755_),
    .A2(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3967_ (.I(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3968_ (.I(_0959_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3969_ (.A1(\mod.registers.r6[6] ),
    .A2(_0684_),
    .B1(_0710_),
    .B2(\mod.registers.r15[6] ),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3970_ (.A1(\mod.registers.r5[6] ),
    .A2(_0896_),
    .B1(_0575_),
    .B2(\mod.registers.r9[6] ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3971_ (.A1(\mod.registers.r11[6] ),
    .A2(_3166_),
    .B1(_0578_),
    .B2(\mod.registers.r10[6] ),
    .C1(\mod.registers.r2[6] ),
    .C2(_0922_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3972_ (.A1(_0967_),
    .A2(_0968_),
    .A3(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3973_ (.I(_3130_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3974_ (.A1(_0476_),
    .A2(_0971_),
    .A3(\mod.registers.r8[6] ),
    .A4(_0581_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3975_ (.A1(_3141_),
    .A2(_3180_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3976_ (.A1(_3173_),
    .A2(_0580_),
    .A3(\mod.registers.r1[6] ),
    .A4(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3977_ (.A1(_0972_),
    .A2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3978_ (.I(\mod.registers.r14[6] ),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(_0585_),
    .A2(_0586_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3980_ (.I(\mod.registers.r7[6] ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3981_ (.A1(_3181_),
    .A2(_0580_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3982_ (.A1(_0885_),
    .A2(_3180_),
    .A3(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3983_ (.A1(_0976_),
    .A2(_0977_),
    .A3(_3179_),
    .B1(_0978_),
    .B2(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3984_ (.I(_3173_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3985_ (.A1(_0982_),
    .A2(_0445_),
    .A3(\mod.registers.r13[6] ),
    .A4(_0583_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3986_ (.A1(\mod.registers.r12[6] ),
    .A2(_0581_),
    .A3(_0583_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3987_ (.A1(_0983_),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3988_ (.A1(\mod.registers.r3[6] ),
    .A2(_0979_),
    .A3(_0973_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3989_ (.A1(_0885_),
    .A2(_0697_),
    .A3(\mod.registers.r4[6] ),
    .A4(_0581_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3990_ (.A1(_0986_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3991_ (.A1(_0975_),
    .A2(_0981_),
    .A3(_0985_),
    .A4(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3992_ (.A1(_0442_),
    .A2(_0970_),
    .A3(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3993_ (.I(_0886_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3994_ (.I0(_0596_),
    .I1(\mod.funct3[1] ),
    .S(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3995_ (.A1(_0966_),
    .A2(_0990_),
    .B1(_0992_),
    .B2(_3222_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3996_ (.A1(_0766_),
    .A2(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3997_ (.A1(_0965_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3998_ (.A1(_0774_),
    .A2(_0779_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3999_ (.A1(\mod.pc_2[5] ),
    .A2(_0594_),
    .B(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4000_ (.A1(\mod.registers.r5[5] ),
    .A2(_0896_),
    .B1(_3172_),
    .B2(\mod.registers.r13[5] ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4001_ (.A1(\mod.registers.r7[5] ),
    .A2(_3134_),
    .B1(_3148_),
    .B2(\mod.registers.r1[5] ),
    .C1(_3166_),
    .C2(\mod.registers.r11[5] ),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4002_ (.A1(\mod.registers.r2[5] ),
    .A2(_0922_),
    .B1(_3139_),
    .B2(\mod.registers.r3[5] ),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4003_ (.A1(_0998_),
    .A2(_0999_),
    .A3(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4004_ (.A1(\mod.registers.r4[5] ),
    .A2(_0565_),
    .B1(_0686_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4005_ (.A1(\mod.registers.r8[5] ),
    .A2(_3168_),
    .B1(_0711_),
    .B2(\mod.registers.r9[5] ),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4006_ (.A1(\mod.registers.r6[5] ),
    .A2(_0572_),
    .B1(_0716_),
    .B2(\mod.registers.r12[5] ),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4007_ (.A1(\mod.registers.r14[5] ),
    .A2(_3176_),
    .B1(_0710_),
    .B2(\mod.registers.r15[5] ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4008_ (.A1(_1003_),
    .A2(_1004_),
    .A3(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4009_ (.A1(_0696_),
    .A2(_1001_),
    .A3(_1002_),
    .A4(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4010_ (.I0(_0889_),
    .I1(\mod.funct7[1] ),
    .S(_0595_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4011_ (.A1(_0696_),
    .A2(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4012_ (.A1(_3221_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4013_ (.I0(_0448_),
    .I1(\mod.funct3[0] ),
    .S(_0886_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4014_ (.A1(_1007_),
    .A2(_1010_),
    .B1(_1011_),
    .B2(_0535_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4015_ (.A1(_0997_),
    .A2(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4016_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4017_ (.A1(_0794_),
    .A2(_0723_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_0781_),
    .A2(_1012_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4019_ (.A1(_1014_),
    .A2(_1015_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4020_ (.I(_0993_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4021_ (.A1(_0767_),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4022_ (.A1(_0755_),
    .A2(_0960_),
    .A3(_0962_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4023_ (.A1(_0965_),
    .A2(_1019_),
    .B(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4024_ (.A1(_0995_),
    .A2(_1017_),
    .B(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4025_ (.A1(_0701_),
    .A2(_0825_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4026_ (.I(\mod.pc_2[3] ),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4027_ (.A1(_0800_),
    .A2(_0801_),
    .A3(_0802_),
    .A4(_0803_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4028_ (.A1(_0805_),
    .A2(_0806_),
    .A3(_0807_),
    .A4(_0809_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4029_ (.A1(_1024_),
    .A2(_3203_),
    .B1(_1025_),
    .B2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4030_ (.A1(_0535_),
    .A2(_0479_),
    .A3(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4031_ (.I(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4032_ (.A1(_0467_),
    .A2(_0475_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4033_ (.A1(_0706_),
    .A2(_0477_),
    .B1(_1030_),
    .B2(_3199_),
    .C(_0811_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4034_ (.A1(_1029_),
    .A2(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4035_ (.A1(_0480_),
    .A2(_0811_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4036_ (.A1(_1023_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4037_ (.I(_0599_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4038_ (.A1(_1035_),
    .A2(_0842_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4039_ (.A1(_0593_),
    .A2(_0598_),
    .B(_0841_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4040_ (.I(\mod.pc_2[1] ),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4041_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0833_),
    .A4(_0834_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4042_ (.A1(_0836_),
    .A2(_0837_),
    .A3(_0838_),
    .A4(_0839_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4043_ (.A1(_1038_),
    .A2(_0453_),
    .B1(_1039_),
    .B2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4044_ (.A1(_3223_),
    .A2(_0844_),
    .A3(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4045_ (.A1(_1037_),
    .A2(_1042_),
    .B1(_0440_),
    .B2(_0562_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4046_ (.A1(_0814_),
    .A2(_0815_),
    .A3(_0816_),
    .A4(_0817_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4047_ (.A1(_0819_),
    .A2(_0820_),
    .A3(_0821_),
    .A4(_0822_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4048_ (.A1(\mod.pc_2[2] ),
    .A2(_0594_),
    .B1(_1044_),
    .B2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4049_ (.A1(_3226_),
    .A2(_0700_),
    .A3(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4050_ (.I(_0564_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4051_ (.A1(_0683_),
    .A2(_0695_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4052_ (.I(_0725_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4053_ (.A1(_1048_),
    .A2(_0698_),
    .B1(_1049_),
    .B2(_1050_),
    .C(_0824_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4054_ (.A1(_1047_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4055_ (.A1(_1036_),
    .A2(_1043_),
    .B(_1052_),
    .C(_1032_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4056_ (.A1(_0965_),
    .A2(_0994_),
    .A3(_1013_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4057_ (.A1(_0792_),
    .A2(_0793_),
    .B1(_0722_),
    .B2(_0705_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4058_ (.A1(_3222_),
    .A2(_0792_),
    .A3(_0722_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4059_ (.I(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4060_ (.A1(_1055_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4061_ (.A1(_1034_),
    .A2(_1053_),
    .B(_1054_),
    .C(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4062_ (.A1(\mod.registers.r12[11] ),
    .A2(_0905_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4063_ (.A1(\mod.registers.r7[11] ),
    .A2(_0892_),
    .B1(_0919_),
    .B2(\mod.registers.r15[11] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4064_ (.A1(\mod.registers.r3[11] ),
    .A2(_0899_),
    .B1(_0894_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4065_ (.A1(\mod.registers.r5[11] ),
    .A2(_0897_),
    .B1(_0907_),
    .B2(\mod.registers.r4[11] ),
    .C1(_0909_),
    .C2(\mod.registers.r8[11] ),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4066_ (.A1(_1060_),
    .A2(_1061_),
    .A3(_1062_),
    .A4(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4067_ (.A1(\mod.registers.r14[11] ),
    .A2(_0917_),
    .B1(_0930_),
    .B2(\mod.registers.r9[11] ),
    .C1(\mod.registers.r2[11] ),
    .C2(_0923_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4068_ (.A1(\mod.registers.r11[11] ),
    .A2(_0916_),
    .B1(_0925_),
    .B2(\mod.registers.r1[11] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4069_ (.A1(\mod.registers.r6[11] ),
    .A2(_0902_),
    .B1(_0928_),
    .B2(\mod.registers.r13[11] ),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4070_ (.A1(_1065_),
    .A2(_1066_),
    .A3(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4071_ (.A1(_1048_),
    .A2(_1064_),
    .A3(_1068_),
    .B(_0966_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4072_ (.A1(_0420_),
    .A2(_0887_),
    .B(_0890_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(_0464_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4074_ (.A1(_1069_),
    .A2(_1071_),
    .B(_0630_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4075_ (.A1(_0630_),
    .A2(_1069_),
    .A3(_1071_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4076_ (.A1(_1072_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4077_ (.A1(\mod.registers.r6[10] ),
    .A2(_0684_),
    .B1(_0566_),
    .B2(\mod.registers.r1[10] ),
    .C1(_0689_),
    .C2(\mod.registers.r13[10] ),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4078_ (.A1(\mod.registers.r2[10] ),
    .A2(_0569_),
    .B1(_0575_),
    .B2(\mod.registers.r9[10] ),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4079_ (.A1(\mod.registers.r11[10] ),
    .A2(_0577_),
    .B1(_0690_),
    .B2(\mod.registers.r14[10] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4080_ (.A1(_1075_),
    .A2(_1076_),
    .A3(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4081_ (.A1(\mod.registers.r3[10] ),
    .A2(_0680_),
    .B1(_0686_),
    .B2(\mod.registers.r10[10] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4082_ (.A1(\mod.registers.r12[10] ),
    .A2(_0716_),
    .B1(_0574_),
    .B2(\mod.registers.r8[10] ),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4083_ (.A1(\mod.registers.r7[10] ),
    .A2(_0679_),
    .B1(_0710_),
    .B2(\mod.registers.r15[10] ),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4084_ (.A1(\mod.registers.r5[10] ),
    .A2(_0568_),
    .B1(_0565_),
    .B2(\mod.registers.r4[10] ),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4085_ (.A1(_1079_),
    .A2(_1080_),
    .A3(_1081_),
    .A4(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4086_ (.A1(_0706_),
    .A2(_1078_),
    .A3(_1083_),
    .B(_0966_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4087_ (.A1(_0991_),
    .A2(_1008_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4088_ (.A1(_0616_),
    .A2(_0991_),
    .B(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4089_ (.A1(_0463_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4090_ (.A1(_1084_),
    .A2(_1087_),
    .B(_0649_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4091_ (.I(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4092_ (.A1(_0649_),
    .A2(_1084_),
    .A3(_1087_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4093_ (.A1(_1089_),
    .A2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4094_ (.I(\mod.pc_2[8] ),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4095_ (.A1(_0670_),
    .A2(_0675_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4096_ (.A1(_1092_),
    .A2(_0678_),
    .B(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4097_ (.A1(\mod.registers.r7[8] ),
    .A2(_0892_),
    .B1(_0928_),
    .B2(\mod.registers.r13[8] ),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4098_ (.A1(\mod.registers.r12[8] ),
    .A2(_0904_),
    .B1(_0917_),
    .B2(\mod.registers.r14[8] ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4099_ (.A1(\mod.registers.r5[8] ),
    .A2(_0897_),
    .B1(_0923_),
    .B2(\mod.registers.r2[8] ),
    .C1(_0915_),
    .C2(\mod.registers.r11[8] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4100_ (.A1(_1095_),
    .A2(_1096_),
    .A3(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4101_ (.A1(\mod.registers.r4[8] ),
    .A2(_0907_),
    .B1(_0930_),
    .B2(\mod.registers.r9[8] ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4102_ (.A1(\mod.registers.r3[8] ),
    .A2(_0899_),
    .B1(_0909_),
    .B2(\mod.registers.r8[8] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4103_ (.A1(\mod.registers.r6[8] ),
    .A2(_0902_),
    .B1(_0894_),
    .B2(\mod.registers.r10[8] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4104_ (.A1(\mod.registers.r1[8] ),
    .A2(_0925_),
    .B1(_0919_),
    .B2(\mod.registers.r15[8] ),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4105_ (.A1(_1100_),
    .A2(_1101_),
    .A3(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4106_ (.A1(_0914_),
    .A2(_1098_),
    .A3(_1099_),
    .A4(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4107_ (.I0(_0477_),
    .I1(_0609_),
    .S(_0991_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4108_ (.A1(_0457_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4109_ (.A1(_0935_),
    .A2(_1104_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4110_ (.A1(_1094_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4111_ (.A1(_1094_),
    .A2(_1107_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4112_ (.A1(_1108_),
    .A2(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4113_ (.I(_0661_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4114_ (.A1(\mod.registers.r13[9] ),
    .A2(_0928_),
    .B1(_0925_),
    .B2(\mod.registers.r1[9] ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4115_ (.A1(\mod.registers.r7[9] ),
    .A2(_0892_),
    .B1(_0923_),
    .B2(\mod.registers.r2[9] ),
    .C1(_0915_),
    .C2(\mod.registers.r11[9] ),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4116_ (.A1(\mod.registers.r4[9] ),
    .A2(_0907_),
    .B1(_0917_),
    .B2(\mod.registers.r14[9] ),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4117_ (.A1(_1112_),
    .A2(_1113_),
    .A3(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4118_ (.A1(\mod.registers.r10[9] ),
    .A2(_0894_),
    .B1(_0930_),
    .B2(\mod.registers.r9[9] ),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4119_ (.A1(\mod.registers.r5[9] ),
    .A2(_0897_),
    .B1(_0899_),
    .B2(\mod.registers.r3[9] ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4120_ (.A1(\mod.registers.r6[9] ),
    .A2(_0902_),
    .B1(_0909_),
    .B2(\mod.registers.r8[9] ),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4121_ (.A1(\mod.registers.r12[9] ),
    .A2(_0904_),
    .B1(_0919_),
    .B2(\mod.registers.r15[9] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4122_ (.A1(_1116_),
    .A2(_1117_),
    .A3(_1118_),
    .A4(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4123_ (.A1(_0564_),
    .A2(_1115_),
    .A3(_1120_),
    .B(_0966_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4124_ (.I0(_0720_),
    .I1(_0608_),
    .S(_0887_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4125_ (.A1(_0457_),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4126_ (.A1(_1121_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4127_ (.A1(_1111_),
    .A2(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4128_ (.A1(_1074_),
    .A2(_1091_),
    .A3(_1110_),
    .A4(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4129_ (.A1(_1022_),
    .A2(_1059_),
    .B(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4130_ (.A1(_1088_),
    .A2(_1090_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4131_ (.A1(_0676_),
    .A2(_1107_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4132_ (.A1(_1111_),
    .A2(_1121_),
    .A3(_1123_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4133_ (.A1(_1125_),
    .A2(_1129_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4134_ (.I(_0649_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4135_ (.A1(_1132_),
    .A2(_1084_),
    .A3(_1087_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4136_ (.A1(_1128_),
    .A2(_1131_),
    .B(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4137_ (.I(_0631_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4138_ (.A1(_1135_),
    .A2(_1069_),
    .A3(_1071_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4139_ (.A1(_1074_),
    .A2(_1134_),
    .B(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4140_ (.I(\mod.pc_2[12] ),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4141_ (.A1(_0554_),
    .A2(_0555_),
    .A3(_0556_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4142_ (.A1(_0547_),
    .A2(_0550_),
    .A3(_0552_),
    .A4(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4143_ (.A1(_1138_),
    .A2(_3223_),
    .B1(_0559_),
    .B2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4144_ (.I(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4145_ (.A1(\mod.registers.r4[12] ),
    .A2(_0908_),
    .B1(_0918_),
    .B2(\mod.registers.r14[12] ),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4146_ (.A1(\mod.registers.r7[12] ),
    .A2(_0893_),
    .B1(_0926_),
    .B2(\mod.registers.r1[12] ),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4147_ (.A1(\mod.registers.r6[12] ),
    .A2(_0903_),
    .B1(_0900_),
    .B2(\mod.registers.r3[12] ),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4148_ (.A1(\mod.registers.r10[12] ),
    .A2(_0895_),
    .B1(_0931_),
    .B2(\mod.registers.r9[12] ),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4149_ (.A1(_1143_),
    .A2(_1144_),
    .A3(_1145_),
    .A4(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4150_ (.A1(\mod.registers.r12[12] ),
    .A2(_0904_),
    .B1(_0924_),
    .B2(\mod.registers.r2[12] ),
    .C1(_0915_),
    .C2(\mod.registers.r11[12] ),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4151_ (.A1(\mod.registers.r13[12] ),
    .A2(_0929_),
    .B1(_0910_),
    .B2(\mod.registers.r8[12] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4152_ (.A1(\mod.registers.r5[12] ),
    .A2(_0898_),
    .B1(_0920_),
    .B2(\mod.registers.r15[12] ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4153_ (.A1(_1148_),
    .A2(_1149_),
    .A3(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4154_ (.A1(_1147_),
    .A2(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4155_ (.A1(_1048_),
    .A2(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4156_ (.A1(_0586_),
    .A2(_1050_),
    .A3(_0934_),
    .B1(_0935_),
    .B2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4157_ (.A1(_1142_),
    .A2(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4158_ (.I(_1154_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4159_ (.A1(_0561_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_1155_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4161_ (.A1(_1127_),
    .A2(_1137_),
    .B(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4162_ (.A1(\mod.registers.r12[13] ),
    .A2(_0905_),
    .B1(_0924_),
    .B2(\mod.registers.r2[13] ),
    .C1(_0900_),
    .C2(\mod.registers.r3[13] ),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4163_ (.A1(\mod.registers.r8[13] ),
    .A2(_0910_),
    .B1(_0920_),
    .B2(\mod.registers.r15[13] ),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4164_ (.A1(\mod.registers.r6[13] ),
    .A2(_0903_),
    .B1(_0898_),
    .B2(\mod.registers.r5[13] ),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4165_ (.A1(\mod.registers.r4[13] ),
    .A2(_0908_),
    .B1(_0895_),
    .B2(\mod.registers.r10[13] ),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4166_ (.A1(\mod.registers.r11[13] ),
    .A2(_0916_),
    .B1(_0926_),
    .B2(\mod.registers.r1[13] ),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4167_ (.A1(\mod.registers.r13[13] ),
    .A2(_0929_),
    .B1(_0931_),
    .B2(\mod.registers.r9[13] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4168_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4169_ (.A1(\mod.registers.r7[13] ),
    .A2(_0893_),
    .B1(_0918_),
    .B2(\mod.registers.r14[13] ),
    .C(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4170_ (.A1(_1160_),
    .A2(_1161_),
    .A3(_1162_),
    .A4(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4171_ (.A1(_1048_),
    .A2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4172_ (.A1(_0982_),
    .A2(_1050_),
    .A3(_0934_),
    .B1(_0935_),
    .B2(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4173_ (.I(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4174_ (.I(_1142_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_1172_),
    .A2(_1156_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4176_ (.A1(_0544_),
    .A2(_1171_),
    .B(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4177_ (.I(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4178_ (.I(_3205_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4179_ (.I(_0889_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4180_ (.A1(_0971_),
    .A2(_0888_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4181_ (.A1(_1177_),
    .A2(_0888_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4182_ (.I(_0531_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4183_ (.A1(\mod.registers.r4[14] ),
    .A2(_0908_),
    .B1(_0926_),
    .B2(\mod.registers.r1[14] ),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4184_ (.A1(\mod.registers.r5[14] ),
    .A2(_0898_),
    .B1(_0924_),
    .B2(\mod.registers.r2[14] ),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4185_ (.A1(\mod.registers.r7[14] ),
    .A2(_0893_),
    .B1(_0929_),
    .B2(\mod.registers.r13[14] ),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4186_ (.A1(\mod.registers.r10[14] ),
    .A2(_0895_),
    .B1(_0931_),
    .B2(\mod.registers.r9[14] ),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4187_ (.A1(_1181_),
    .A2(_1182_),
    .A3(_1183_),
    .A4(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4188_ (.A1(\mod.registers.r12[14] ),
    .A2(_0905_),
    .B1(_0900_),
    .B2(\mod.registers.r3[14] ),
    .C1(_0910_),
    .C2(\mod.registers.r8[14] ),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4189_ (.A1(\mod.registers.r11[14] ),
    .A2(_0916_),
    .B1(_0918_),
    .B2(\mod.registers.r14[14] ),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4190_ (.A1(\mod.registers.r6[14] ),
    .A2(_0903_),
    .B1(_0920_),
    .B2(\mod.registers.r15[14] ),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4191_ (.A1(_1186_),
    .A2(_1187_),
    .A3(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4192_ (.A1(_1185_),
    .A2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4193_ (.A1(_0914_),
    .A2(_1190_),
    .B(_0958_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4194_ (.A1(_1176_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4195_ (.A1(_1176_),
    .A2(_1179_),
    .B(_1180_),
    .C(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4196_ (.A1(_0525_),
    .A2(_0530_),
    .B(_1176_),
    .C(_1191_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4197_ (.A1(_1193_),
    .A2(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_0544_),
    .A2(_1171_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4199_ (.I(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4200_ (.A1(_1159_),
    .A2(_1175_),
    .B(_1195_),
    .C(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4201_ (.A1(_1191_),
    .A2(_1180_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4202_ (.A1(_0943_),
    .A2(_1198_),
    .A3(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4203_ (.A1(_1198_),
    .A2(_1199_),
    .B(_0943_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4204_ (.A1(_0728_),
    .A2(_0731_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4205_ (.I(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4206_ (.I(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4208_ (.A1(_1200_),
    .A2(_1201_),
    .B(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4209_ (.I(_0732_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4210_ (.I(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4211_ (.I(\mod.pc_2[13] ),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4212_ (.A1(_1209_),
    .A2(_0464_),
    .B1(_0537_),
    .B2(_0542_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4213_ (.I(_1210_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4214_ (.A1(_1211_),
    .A2(_1171_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4215_ (.A1(_1211_),
    .A2(_1171_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4216_ (.A1(_1155_),
    .A2(_1212_),
    .B(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4217_ (.A1(_0965_),
    .A2(_0994_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4218_ (.I(_1047_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4219_ (.A1(_0480_),
    .A2(_1027_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4220_ (.A1(_0593_),
    .A2(_0598_),
    .A3(_0841_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4221_ (.A1(_1218_),
    .A2(_0867_),
    .B(_1037_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4222_ (.A1(_1047_),
    .A2(_1051_),
    .A3(_1029_),
    .A4(_1031_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4223_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_1219_),
    .B2(_1220_),
    .C(_1029_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4224_ (.A1(_1055_),
    .A2(_1056_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4225_ (.A1(_1014_),
    .A2(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4226_ (.I(_0964_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4227_ (.I(_0994_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4228_ (.I(_0997_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4229_ (.I(_1012_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4230_ (.A1(_1226_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4231_ (.A1(_1226_),
    .A2(_1227_),
    .B(_1057_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4232_ (.A1(_1224_),
    .A2(_1225_),
    .A3(_1228_),
    .A4(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4233_ (.A1(_1215_),
    .A2(_1221_),
    .A3(_1223_),
    .B(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4234_ (.I(_0755_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4235_ (.A1(_1232_),
    .A2(_0963_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4236_ (.I(_0766_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4237_ (.A1(_1234_),
    .A2(_1018_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4238_ (.A1(_1232_),
    .A2(_0963_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4239_ (.A1(_1233_),
    .A2(_1235_),
    .B(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4240_ (.I(_1128_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4241_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4242_ (.I(_1111_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4243_ (.A1(_1240_),
    .A2(_1124_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4244_ (.A1(_0662_),
    .A2(_1121_),
    .A3(_1123_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4245_ (.A1(_1241_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4246_ (.A1(_1238_),
    .A2(_1239_),
    .A3(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4247_ (.I(_1074_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4248_ (.A1(_1231_),
    .A2(_1237_),
    .B(_1244_),
    .C(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4249_ (.I(_1089_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4250_ (.A1(_1094_),
    .A2(_1107_),
    .A3(_1242_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4251_ (.A1(_1241_),
    .A2(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4252_ (.A1(_1247_),
    .A2(_1249_),
    .B(_1090_),
    .C(_1073_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4253_ (.A1(_1072_),
    .A2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4254_ (.A1(_0544_),
    .A2(_1170_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4255_ (.A1(_1246_),
    .A2(_1251_),
    .B(_1158_),
    .C(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4256_ (.A1(_1214_),
    .A2(_1253_),
    .B(_1195_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4257_ (.A1(_0942_),
    .A2(_1194_),
    .A3(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4258_ (.A1(_1194_),
    .A2(_1254_),
    .B(_0942_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4259_ (.A1(_1208_),
    .A2(_1255_),
    .A3(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4260_ (.I(_0875_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4261_ (.I(_0861_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4262_ (.I(_0866_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4263_ (.I(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4264_ (.A1(_0941_),
    .A2(_1261_),
    .B(_0947_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4265_ (.A1(_0940_),
    .A2(_1259_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4266_ (.I(_0856_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4267_ (.I(_0828_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4268_ (.I(_1035_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4269_ (.I(_0826_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4270_ (.A1(_1266_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4271_ (.A1(_1265_),
    .A2(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4272_ (.I(_0482_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4273_ (.I(_0458_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4274_ (.A1(_0939_),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4275_ (.I(_0847_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4276_ (.I(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4277_ (.A1(_1270_),
    .A2(_1272_),
    .A3(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4278_ (.A1(_0853_),
    .A2(_0722_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4279_ (.A1(_1276_),
    .A2(_0735_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4280_ (.A1(_1277_),
    .A2(_0733_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4281_ (.I(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4282_ (.A1(_0733_),
    .A2(_1269_),
    .B(_1275_),
    .C(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4283_ (.I(_0737_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(_0701_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4285_ (.I(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4286_ (.I(_0846_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4288_ (.I(_1041_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4289_ (.I(_0796_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4290_ (.A1(_1286_),
    .A2(_1287_),
    .B(_0452_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4291_ (.A1(_1285_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4292_ (.I(_1035_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4293_ (.A1(_0812_),
    .A2(_1287_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4294_ (.A1(_1267_),
    .A2(_1046_),
    .B(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_1290_),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(_1289_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4297_ (.I(_0701_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4299_ (.A1(\mod.pc_2[7] ),
    .A2(_1176_),
    .B1(_0745_),
    .B2(_0753_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4300_ (.I(_0459_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4301_ (.I(_1298_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4302_ (.I(_3223_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4303_ (.I(_0451_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4304_ (.A1(_1300_),
    .A2(_1234_),
    .A3(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4305_ (.A1(_1297_),
    .A2(_1299_),
    .B(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4306_ (.I(_0845_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4307_ (.A1(_1300_),
    .A2(_1301_),
    .B(_0781_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4308_ (.I(_0459_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4309_ (.A1(_0795_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4310_ (.A1(_1304_),
    .A2(_1305_),
    .A3(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4311_ (.A1(_1285_),
    .A2(_1303_),
    .B(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4312_ (.A1(_1296_),
    .A2(_1309_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4313_ (.A1(_1283_),
    .A2(_1294_),
    .B(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_0828_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4315_ (.I(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(_1094_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4317_ (.A1(_1306_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4318_ (.A1(_1306_),
    .A2(_0662_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4319_ (.I(_0797_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4320_ (.I0(_0631_),
    .I1(_0650_),
    .S(_1298_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4321_ (.A1(_1317_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4322_ (.A1(_1290_),
    .A2(_1316_),
    .B(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4323_ (.A1(_1300_),
    .A2(_1301_),
    .B(_1210_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4324_ (.A1(_1172_),
    .A2(_1299_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4325_ (.A1(_1321_),
    .A2(_1322_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4326_ (.I(_0829_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4327_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4328_ (.A1(_0853_),
    .A2(_0531_),
    .A3(_0451_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4329_ (.A1(_0883_),
    .A2(_1267_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4330_ (.A1(_1326_),
    .A2(_1327_),
    .A3(_1273_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4331_ (.A1(_1313_),
    .A2(_1320_),
    .B1(_1323_),
    .B2(_1325_),
    .C(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4332_ (.A1(_1281_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4333_ (.A1(_1281_),
    .A2(_1311_),
    .B(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4334_ (.A1(_0945_),
    .A2(_0855_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4335_ (.A1(_1264_),
    .A2(_1280_),
    .B1(_1331_),
    .B2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4336_ (.A1(_0942_),
    .A2(_1258_),
    .B(_1263_),
    .C(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4337_ (.A1(_1200_),
    .A2(_1201_),
    .B(_3210_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4338_ (.A1(_0948_),
    .A2(_1206_),
    .A3(_1257_),
    .B1(_1334_),
    .B2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4339_ (.I(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4340_ (.A1(_0884_),
    .A2(_0937_),
    .B1(_0943_),
    .B2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4341_ (.A1(_0874_),
    .A2(_1337_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4342_ (.A1(_3192_),
    .A2(_3207_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4343_ (.I(_1340_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4345_ (.A1(_0874_),
    .A2(_1338_),
    .B(_1339_),
    .C(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4346_ (.A1(_0880_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4347_ (.I(\mod.valid2 ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4348_ (.I(_1345_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4349_ (.I(_0945_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4350_ (.I(_3193_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4351_ (.A1(_1347_),
    .A2(_1348_),
    .A3(_1338_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(_0865_),
    .A2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4353_ (.A1(_3212_),
    .A2(_1338_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4354_ (.I(_1158_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4355_ (.A1(_1127_),
    .A2(_1137_),
    .A3(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(_1202_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4357_ (.I(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4358_ (.A1(_1355_),
    .A2(_0947_),
    .B(_3209_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4359_ (.A1(_1159_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4360_ (.A1(_1353_),
    .A2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4361_ (.I(_1296_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4362_ (.A1(_1306_),
    .A2(_1314_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4363_ (.A1(_1297_),
    .A2(_1299_),
    .B(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4364_ (.A1(_1234_),
    .A2(_0862_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4365_ (.A1(_1226_),
    .A2(_1271_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4366_ (.A1(_1362_),
    .A2(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4367_ (.I0(_1361_),
    .I1(_1364_),
    .S(_1304_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4368_ (.I(_1271_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4369_ (.A1(_1172_),
    .A2(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4370_ (.A1(_1366_),
    .A2(_0631_),
    .B(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4371_ (.I(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4372_ (.I(_0863_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4373_ (.A1(_0863_),
    .A2(_0650_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4374_ (.A1(_1370_),
    .A2(_1240_),
    .B(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4375_ (.I(_0481_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4376_ (.A1(_1373_),
    .A2(_1332_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4377_ (.I(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4378_ (.A1(_1274_),
    .A2(_1369_),
    .B1(_1372_),
    .B2(_1325_),
    .C(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4379_ (.A1(_1359_),
    .A2(_1365_),
    .B(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4380_ (.I(_1264_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4381_ (.I(_0735_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4383_ (.I(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4384_ (.A1(_0882_),
    .A2(_0702_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4385_ (.I(_1276_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4386_ (.A1(_1383_),
    .A2(_1354_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4387_ (.A1(_1265_),
    .A2(_0601_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4388_ (.A1(_1382_),
    .A2(_1384_),
    .B(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(_1279_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4390_ (.A1(_1381_),
    .A2(_1386_),
    .B(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4391_ (.I(_1282_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4392_ (.A1(_0792_),
    .A2(_0793_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4393_ (.I0(_1390_),
    .I1(_1027_),
    .I2(_1046_),
    .I3(_1286_),
    .S0(_1271_),
    .S1(_1284_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4394_ (.A1(_1317_),
    .A2(_0460_),
    .B(_1295_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4395_ (.A1(_1389_),
    .A2(_1391_),
    .B(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4396_ (.I(_0871_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4397_ (.A1(_0482_),
    .A2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4398_ (.I(_0875_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4399_ (.A1(_3207_),
    .A2(_0859_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4400_ (.A1(_1155_),
    .A2(_1260_),
    .B(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4401_ (.A1(_1157_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4402_ (.A1(_1352_),
    .A2(_1396_),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4403_ (.A1(_1378_),
    .A2(_1388_),
    .B1(_1393_),
    .B2(_1395_),
    .C(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4404_ (.A1(_1377_),
    .A2(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4405_ (.A1(_1246_),
    .A2(_1251_),
    .B(_1352_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4406_ (.A1(_1352_),
    .A2(_1246_),
    .A3(_1251_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4407_ (.A1(_1208_),
    .A2(_0948_),
    .A3(_1403_),
    .A4(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4408_ (.A1(_1358_),
    .A2(_1402_),
    .A3(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_1125_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4410_ (.I(_1129_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_1110_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4412_ (.A1(_1022_),
    .A2(_1059_),
    .B(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4413_ (.A1(_1408_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4414_ (.A1(_1407_),
    .A2(_1411_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4415_ (.I(_1108_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4416_ (.A1(_1231_),
    .A2(_1237_),
    .B(_1409_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4417_ (.A1(_1413_),
    .A2(_1414_),
    .B(_1407_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4418_ (.A1(_1413_),
    .A2(_1407_),
    .A3(_1414_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(_1355_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4420_ (.I(_0869_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4421_ (.A1(_1205_),
    .A2(_1412_),
    .B1(_1415_),
    .B2(_1417_),
    .C(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4422_ (.I(_1341_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(_1420_),
    .A2(_1412_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4424_ (.I(_1035_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4425_ (.A1(_1422_),
    .A2(_1305_),
    .A3(_1307_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4426_ (.A1(_1317_),
    .A2(_1292_),
    .B(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4427_ (.I0(_1303_),
    .I1(_1316_),
    .S(_1290_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4428_ (.A1(_1283_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4429_ (.I(_1373_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4430_ (.A1(_1359_),
    .A2(_1424_),
    .B(_1426_),
    .C(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4431_ (.A1(_1288_),
    .A2(_1274_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4432_ (.A1(_1381_),
    .A2(_1429_),
    .B(_1394_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4433_ (.A1(_1241_),
    .A2(_1261_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4434_ (.A1(_1242_),
    .A2(_1259_),
    .B1(_1428_),
    .B2(_1430_),
    .C(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4435_ (.A1(_1348_),
    .A2(_0944_),
    .A3(_0881_),
    .A4(_0859_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4436_ (.I(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4437_ (.A1(_0882_),
    .A2(_0797_),
    .A3(_0702_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_1366_),
    .A2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(_1207_),
    .A2(_1277_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4440_ (.I(_0739_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_1438_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4442_ (.A1(_1266_),
    .A2(_1326_),
    .A3(_1321_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4443_ (.A1(_1422_),
    .A2(_1272_),
    .B(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4444_ (.I0(_1141_),
    .I1(_1135_),
    .I2(_1132_),
    .I3(_1240_),
    .S0(_0796_),
    .S1(_0600_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4445_ (.A1(_0739_),
    .A2(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4446_ (.A1(_1439_),
    .A2(_1441_),
    .B(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4447_ (.A1(_1427_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4448_ (.A1(_1436_),
    .A2(_1437_),
    .B(_1445_),
    .C(_1387_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4449_ (.A1(_1407_),
    .A2(_1434_),
    .B1(_1446_),
    .B2(_1378_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4450_ (.A1(_1419_),
    .A2(_1421_),
    .A3(_1432_),
    .A4(_1447_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4451_ (.A1(_1409_),
    .A2(_1231_),
    .A3(_1237_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4452_ (.A1(_1449_),
    .A2(_1414_),
    .B(_1207_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4453_ (.A1(_1022_),
    .A2(_1059_),
    .B(_1239_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4454_ (.I(_1224_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4455_ (.A1(_0780_),
    .A2(_1012_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4456_ (.I(_1453_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4457_ (.A1(_1390_),
    .A2(_1383_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4458_ (.A1(_0781_),
    .A2(_1227_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4459_ (.A1(_1454_),
    .A2(_1455_),
    .B(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4460_ (.A1(_1224_),
    .A2(_1225_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4461_ (.A1(_1452_),
    .A2(_1019_),
    .B1(_1457_),
    .B2(_1458_),
    .C(_1020_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4462_ (.A1(_0738_),
    .A2(_1046_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4463_ (.A1(_1028_),
    .A2(_1031_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4464_ (.I(_1461_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4465_ (.A1(_0735_),
    .A2(_1027_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4466_ (.A1(_1460_),
    .A2(_1462_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4467_ (.A1(_0845_),
    .A2(_1286_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4468_ (.A1(_0705_),
    .A2(_0844_),
    .B(_1286_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4469_ (.A1(_1466_),
    .A2(_1218_),
    .B(_0452_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4470_ (.A1(_1047_),
    .A2(_1051_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4471_ (.A1(_1465_),
    .A2(_1467_),
    .B(_1468_),
    .C(_1461_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4472_ (.A1(_1224_),
    .A2(_1225_),
    .A3(_1014_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4473_ (.A1(_1464_),
    .A2(_1469_),
    .B(_1470_),
    .C(_1222_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4474_ (.A1(_1459_),
    .A2(_1471_),
    .A3(_1409_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4475_ (.A1(_1204_),
    .A2(_1451_),
    .A3(_1472_),
    .B(_1418_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4476_ (.A1(_1451_),
    .A2(_1472_),
    .B(_1341_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4477_ (.A1(_0737_),
    .A2(_0703_),
    .B(_1279_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_0857_),
    .A2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4479_ (.I(_0739_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_1477_),
    .A2(_1391_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4481_ (.I(_0872_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4482_ (.A1(_1313_),
    .A2(_1365_),
    .B(_1478_),
    .C(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4483_ (.A1(_1413_),
    .A2(_1433_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4484_ (.A1(_1413_),
    .A2(_0866_),
    .B(_1481_),
    .C(_1397_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4485_ (.A1(_1109_),
    .A2(_1482_),
    .B1(_0873_),
    .B2(_1395_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4486_ (.A1(_1476_),
    .A2(_1480_),
    .A3(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4487_ (.A1(_1450_),
    .A2(_1473_),
    .B(_1474_),
    .C(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4488_ (.I(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4489_ (.A1(_1464_),
    .A2(_1469_),
    .B(_1222_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4490_ (.A1(_1487_),
    .A2(_1455_),
    .B(_1453_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4491_ (.I(_1058_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4492_ (.A1(_1034_),
    .A2(_1053_),
    .B(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4493_ (.A1(_1014_),
    .A2(_1490_),
    .A3(_1015_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4494_ (.A1(_1488_),
    .A2(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4495_ (.A1(_1489_),
    .A2(_1221_),
    .B(_1057_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4496_ (.A1(_1454_),
    .A2(_1493_),
    .B(_1204_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4497_ (.A1(_1454_),
    .A2(_1493_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4498_ (.A1(_1207_),
    .A2(_1492_),
    .B(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4499_ (.A1(_1284_),
    .A2(_1282_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4500_ (.A1(_1477_),
    .A2(_1424_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4501_ (.A1(_1288_),
    .A2(_1497_),
    .B(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4502_ (.A1(_0865_),
    .A2(_3207_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4504_ (.A1(_1226_),
    .A2(_1227_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4505_ (.A1(_1228_),
    .A2(_1259_),
    .B1(_1501_),
    .B2(_1502_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4506_ (.A1(_1454_),
    .A2(_1258_),
    .B1(_1499_),
    .B2(_1375_),
    .C(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4507_ (.A1(_0938_),
    .A2(_1383_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4508_ (.A1(_1266_),
    .A2(_0702_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4509_ (.A1(_0884_),
    .A2(_0723_),
    .A3(_1379_),
    .A4(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4510_ (.A1(_1383_),
    .A2(_0736_),
    .B(_0732_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4511_ (.A1(_1505_),
    .A2(_1507_),
    .B(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4512_ (.A1(_0863_),
    .A2(_1296_),
    .A3(_1505_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4513_ (.A1(_1477_),
    .A2(_1441_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4514_ (.I0(_1232_),
    .I1(_1314_),
    .S(_1298_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4515_ (.A1(_1266_),
    .A2(_1305_),
    .A3(_1302_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4516_ (.A1(_1290_),
    .A2(_1512_),
    .B(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4517_ (.A1(_1389_),
    .A2(_1442_),
    .B(_0481_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4518_ (.A1(_1389_),
    .A2(_1514_),
    .B(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4519_ (.A1(_1509_),
    .A2(_1510_),
    .B1(_1511_),
    .B2(_1281_),
    .C(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4520_ (.I(_0852_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4521_ (.A1(_0945_),
    .A2(_1518_),
    .A3(_0854_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4522_ (.I(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4523_ (.A1(_3209_),
    .A2(_1492_),
    .B1(_1517_),
    .B2(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4524_ (.A1(_1418_),
    .A2(_1496_),
    .B(_1504_),
    .C(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4525_ (.A1(_1055_),
    .A2(_0861_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4526_ (.A1(_1489_),
    .A2(_1396_),
    .B1(_1260_),
    .B2(_1057_),
    .C(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4527_ (.A1(_1312_),
    .A2(_0798_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4528_ (.A1(_1438_),
    .A2(_0677_),
    .B(_1379_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_0736_),
    .A2(_1382_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4530_ (.A1(_1505_),
    .A2(_1527_),
    .B(_1508_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4531_ (.A1(_1380_),
    .A2(_1385_),
    .B1(_1525_),
    .B2(_1526_),
    .C(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4532_ (.A1(_1479_),
    .A2(_1393_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4533_ (.A1(_1520_),
    .A2(_1529_),
    .B(_1530_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4534_ (.A1(_1222_),
    .A2(_1464_),
    .A3(_1469_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4535_ (.A1(_1490_),
    .A2(_1532_),
    .B(_1354_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4536_ (.A1(_1489_),
    .A2(_1221_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4537_ (.A1(_0732_),
    .A2(_1534_),
    .B(_0869_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4538_ (.A1(_1340_),
    .A2(_1490_),
    .A3(_1532_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4539_ (.A1(_1533_),
    .A2(_1535_),
    .B(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4540_ (.A1(_1524_),
    .A2(_1531_),
    .A3(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4541_ (.A1(_1465_),
    .A2(_1467_),
    .B(_1468_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_1539_),
    .A2(_1023_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4543_ (.A1(_1462_),
    .A2(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4544_ (.A1(_1289_),
    .A2(_1293_),
    .B(_1313_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4545_ (.A1(_1029_),
    .A2(_1500_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4546_ (.A1(_1462_),
    .A2(_1396_),
    .B1(_1397_),
    .B2(_1031_),
    .C(_1543_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4547_ (.A1(_1341_),
    .A2(_1541_),
    .B1(_1542_),
    .B2(_1479_),
    .C(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_1506_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4549_ (.I0(_0795_),
    .I1(_0812_),
    .S(_0862_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4550_ (.I0(_1297_),
    .I1(_0676_),
    .I2(_0662_),
    .I3(_0650_),
    .S0(_1298_),
    .S1(_1284_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4551_ (.A1(_1438_),
    .A2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4552_ (.A1(_1305_),
    .A2(_1302_),
    .A3(_1324_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4553_ (.A1(_1546_),
    .A2(_1547_),
    .B(_1549_),
    .C(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4554_ (.A1(_0882_),
    .A2(_0723_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4555_ (.A1(_1268_),
    .A2(_1552_),
    .B(_1528_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4556_ (.I0(_1142_),
    .I1(_1135_),
    .S(_0862_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4557_ (.A1(_1304_),
    .A2(_1326_),
    .A3(_1321_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4558_ (.A1(_1304_),
    .A2(_1554_),
    .B(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4559_ (.A1(_1317_),
    .A2(_1312_),
    .A3(_1272_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4560_ (.A1(_1265_),
    .A2(_1556_),
    .B(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_1380_),
    .A2(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4562_ (.A1(_1281_),
    .A2(_1551_),
    .B(_1553_),
    .C(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4563_ (.A1(_1052_),
    .A2(_1219_),
    .B(_1216_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4564_ (.A1(_1462_),
    .A2(_1561_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4565_ (.I0(_1541_),
    .I1(_1562_),
    .S(_1203_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4566_ (.A1(_1264_),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1418_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4567_ (.A1(_1422_),
    .A2(_1512_),
    .B(_1513_),
    .C(_1312_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4568_ (.I0(_0842_),
    .I1(_0825_),
    .S(_0459_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4569_ (.A1(_1324_),
    .A2(_1547_),
    .B1(_1566_),
    .B2(_0847_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4570_ (.A1(_1565_),
    .A2(_1567_),
    .B(_1379_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4571_ (.A1(_1505_),
    .A2(_1436_),
    .B(_1508_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4572_ (.A1(_1265_),
    .A2(_1441_),
    .B(_1443_),
    .C(_0481_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4573_ (.A1(_1568_),
    .A2(_1569_),
    .A3(_1570_),
    .B(_0857_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4574_ (.A1(_1037_),
    .A2(_1042_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4575_ (.A1(_1572_),
    .A2(_0452_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_1340_),
    .A2(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4577_ (.A1(_1288_),
    .A2(_1273_),
    .A3(_0872_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4578_ (.A1(_1572_),
    .A2(_1433_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4579_ (.A1(_1466_),
    .A2(_0860_),
    .B1(_1500_),
    .B2(_1042_),
    .C(_3216_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4580_ (.A1(_1574_),
    .A2(_1575_),
    .A3(_1576_),
    .A4(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4581_ (.A1(_1299_),
    .A2(_1202_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4582_ (.A1(_1573_),
    .A2(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4583_ (.A1(_1571_),
    .A2(_1578_),
    .B1(_1580_),
    .B2(_3217_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4584_ (.A1(_0795_),
    .A2(_1366_),
    .B(_1363_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4585_ (.I0(_1232_),
    .I1(_0767_),
    .I2(_1240_),
    .I3(_1314_),
    .S0(_0826_),
    .S1(_0846_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4586_ (.A1(_1295_),
    .A2(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4587_ (.A1(_1506_),
    .A2(_0827_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4588_ (.A1(_1324_),
    .A2(_1582_),
    .B(_1584_),
    .C(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4589_ (.A1(_1300_),
    .A2(_0938_),
    .A3(_1301_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4590_ (.A1(_1180_),
    .A2(_1287_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4591_ (.I0(_1211_),
    .I1(_1142_),
    .I2(_1135_),
    .I3(_1132_),
    .S0(_0796_),
    .S1(_0797_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4592_ (.A1(_1588_),
    .A2(_1497_),
    .B1(_1589_),
    .B2(_1282_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4593_ (.A1(_1552_),
    .A2(_1435_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4594_ (.A1(_0482_),
    .A2(_1590_),
    .B1(_1591_),
    .B2(_1508_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4595_ (.A1(_1373_),
    .A2(_1586_),
    .B(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4596_ (.A1(_1036_),
    .A2(_1043_),
    .A3(_1052_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4597_ (.A1(_1539_),
    .A2(_1594_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4598_ (.I0(_0842_),
    .I1(_0825_),
    .S(_0563_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4599_ (.I0(_1596_),
    .I1(_0460_),
    .S(_0846_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4600_ (.A1(_1295_),
    .A2(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4601_ (.A1(_1216_),
    .A2(_0875_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4602_ (.A1(_1216_),
    .A2(_1500_),
    .B(_1599_),
    .C(_0860_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4603_ (.A1(_1051_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4604_ (.A1(_1340_),
    .A2(_1595_),
    .B1(_1598_),
    .B2(_0872_),
    .C(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4605_ (.A1(_1468_),
    .A2(_1219_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_1203_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4607_ (.A1(_1354_),
    .A2(_1595_),
    .B(_1604_),
    .C(_0869_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4608_ (.A1(_1519_),
    .A2(_1593_),
    .B(_1602_),
    .C(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4609_ (.A1(_0879_),
    .A2(_1581_),
    .A3(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4610_ (.A1(_1538_),
    .A2(_1545_),
    .A3(_1564_),
    .A4(_1607_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4611_ (.I(_3217_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_1225_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4613_ (.A1(_1016_),
    .A2(_1488_),
    .B(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4614_ (.A1(_1610_),
    .A2(_1016_),
    .A3(_1488_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4615_ (.A1(_1228_),
    .A2(_1229_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4616_ (.A1(_1221_),
    .A2(_1223_),
    .B(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4617_ (.A1(_1610_),
    .A2(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_1610_),
    .A2(_1614_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_1204_),
    .A2(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4620_ (.A1(_1355_),
    .A2(_1611_),
    .A3(_1612_),
    .B1(_1615_),
    .B2(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4621_ (.A1(_3209_),
    .A2(_1611_),
    .A3(_1612_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_1273_),
    .A2(_1588_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4623_ (.A1(_1389_),
    .A2(_1589_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4624_ (.A1(_1477_),
    .A2(_1583_),
    .B(_1373_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4625_ (.A1(_1270_),
    .A2(_1620_),
    .B1(_1621_),
    .B2(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4626_ (.A1(_1509_),
    .A2(_1623_),
    .B(_1264_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4627_ (.A1(_0812_),
    .A2(_1287_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4628_ (.A1(_1390_),
    .A2(_1267_),
    .B(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4629_ (.I0(_1626_),
    .I1(_1364_),
    .S(_1422_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4630_ (.I0(_1627_),
    .I1(_1597_),
    .S(_1438_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(_1235_),
    .A2(_1434_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(_1397_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4633_ (.A1(_1235_),
    .A2(_1260_),
    .B(_1629_),
    .C(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4634_ (.A1(_1234_),
    .A2(_1018_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4635_ (.A1(_1479_),
    .A2(_1628_),
    .B1(_1631_),
    .B2(_1632_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(_1624_),
    .A2(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4637_ (.A1(_1609_),
    .A2(_1618_),
    .B(_1619_),
    .C(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4638_ (.A1(_1486_),
    .A2(_1522_),
    .A3(_1608_),
    .A4(_1635_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4639_ (.A1(_1406_),
    .A2(_1448_),
    .A3(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4640_ (.I(_1355_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4641_ (.A1(_1408_),
    .A2(_1410_),
    .B(_1243_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4642_ (.A1(_1130_),
    .A2(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4643_ (.A1(_1238_),
    .A2(_1640_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4644_ (.A1(_1231_),
    .A2(_1237_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4645_ (.A1(_1239_),
    .A2(_1243_),
    .A3(_1642_),
    .B(_1249_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4646_ (.A1(_1238_),
    .A2(_1643_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4647_ (.A1(_1205_),
    .A2(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4648_ (.A1(_1638_),
    .A2(_1641_),
    .B(_1645_),
    .C(_1609_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4649_ (.A1(_1208_),
    .A2(_1435_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4650_ (.A1(_1381_),
    .A2(_1590_),
    .B(_1647_),
    .C(_1387_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4651_ (.A1(_1089_),
    .A2(_1501_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4652_ (.A1(_1238_),
    .A2(_1258_),
    .B1(_1630_),
    .B2(_1090_),
    .C(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4653_ (.A1(_1285_),
    .A2(_1361_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4654_ (.A1(_1285_),
    .A2(_1372_),
    .B(_1651_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_1359_),
    .A2(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4656_ (.A1(_1439_),
    .A2(_1627_),
    .B(_1381_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_1427_),
    .A2(_1598_),
    .B(_1332_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4658_ (.A1(_1653_),
    .A2(_1654_),
    .B(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4659_ (.A1(_1378_),
    .A2(_1648_),
    .B(_1650_),
    .C(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_1342_),
    .A2(_1641_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4661_ (.A1(_1646_),
    .A2(_1657_),
    .A3(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_1173_),
    .A2(_1159_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4663_ (.A1(_1660_),
    .A2(_1252_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4664_ (.A1(_1638_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4665_ (.I(_1208_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4666_ (.A1(_1172_),
    .A2(_1154_),
    .B(_1403_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4667_ (.A1(_1252_),
    .A2(_1664_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4668_ (.A1(_1663_),
    .A2(_1665_),
    .B(_1609_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(_1420_),
    .A2(_1661_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4670_ (.A1(_0884_),
    .A2(_1546_),
    .A3(_1384_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4671_ (.A1(_1370_),
    .A2(_1283_),
    .B(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4672_ (.I(_1270_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4673_ (.A1(_1511_),
    .A2(_1669_),
    .B(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_1387_),
    .A2(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4675_ (.A1(_1670_),
    .A2(_1394_),
    .A3(_1499_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4676_ (.A1(_1213_),
    .A2(_1434_),
    .B(_1259_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4677_ (.A1(_1274_),
    .A2(_1323_),
    .B1(_1325_),
    .B2(_1318_),
    .C(_1374_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4678_ (.A1(_1359_),
    .A2(_1425_),
    .B(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4679_ (.A1(_1213_),
    .A2(_1261_),
    .B1(_1674_),
    .B2(_1212_),
    .C(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4680_ (.A1(_1378_),
    .A2(_1672_),
    .B(_1673_),
    .C(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4681_ (.A1(_1662_),
    .A2(_1666_),
    .B(_1667_),
    .C(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4682_ (.I(_1195_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4683_ (.A1(_1159_),
    .A2(_1175_),
    .B(_1197_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4684_ (.A1(_1680_),
    .A2(_1681_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4685_ (.A1(_1211_),
    .A2(_1370_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4686_ (.A1(_1180_),
    .A2(_1370_),
    .B(_1546_),
    .C(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4687_ (.A1(_1325_),
    .A2(_1368_),
    .B1(_1652_),
    .B2(_1439_),
    .C(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(_0884_),
    .A2(_1506_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4689_ (.A1(_0737_),
    .A2(_1620_),
    .B1(_1686_),
    .B2(_1203_),
    .C(_1279_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4690_ (.A1(_0857_),
    .A2(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4691_ (.I(_1194_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4692_ (.A1(_1193_),
    .A2(_0861_),
    .B1(_1501_),
    .B2(_1689_),
    .C(_3217_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4693_ (.A1(_1680_),
    .A2(_1396_),
    .B(_1688_),
    .C(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4694_ (.A1(_1395_),
    .A2(_1628_),
    .B(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4695_ (.A1(_1375_),
    .A2(_1685_),
    .B(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4696_ (.A1(_1420_),
    .A2(_1682_),
    .B(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4697_ (.A1(_1195_),
    .A2(_1214_),
    .A3(_1253_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4698_ (.A1(_1205_),
    .A2(_1254_),
    .A3(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4699_ (.A1(_1663_),
    .A2(_1682_),
    .B(_1696_),
    .C(_0948_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4700_ (.A1(_0767_),
    .A2(_1018_),
    .B(_1611_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4701_ (.A1(_1452_),
    .A2(_1698_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4702_ (.A1(_1638_),
    .A2(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4703_ (.A1(_1235_),
    .A2(_1616_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4704_ (.A1(_1452_),
    .A2(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4705_ (.A1(_1663_),
    .A2(_1702_),
    .B(_1609_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4706_ (.A1(_1296_),
    .A2(_1548_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_1313_),
    .A2(_1556_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4708_ (.A1(_1270_),
    .A2(_1704_),
    .A3(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4709_ (.A1(_1327_),
    .A2(_1546_),
    .B1(_1278_),
    .B2(_1269_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4710_ (.A1(_1380_),
    .A2(_1707_),
    .B(_0734_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4711_ (.A1(_1706_),
    .A2(_1708_),
    .B(_1520_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4712_ (.A1(_1311_),
    .A2(_1375_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4713_ (.A1(_1233_),
    .A2(_1630_),
    .B1(_1261_),
    .B2(_1236_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4714_ (.A1(_1709_),
    .A2(_1710_),
    .A3(_1711_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4715_ (.A1(_1452_),
    .A2(_1434_),
    .B1(_1699_),
    .B2(_1420_),
    .C(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4716_ (.A1(_1694_),
    .A2(_1697_),
    .B1(_1700_),
    .B2(_1703_),
    .C(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4717_ (.A1(_1637_),
    .A2(_1659_),
    .A3(_1679_),
    .A4(_1714_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4718_ (.A1(_1130_),
    .A2(_1639_),
    .B(_1091_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4719_ (.A1(_1133_),
    .A2(_1716_),
    .B(_1245_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4720_ (.A1(_1245_),
    .A2(_1133_),
    .A3(_1716_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4721_ (.A1(_1663_),
    .A2(_1717_),
    .A3(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4722_ (.A1(_1091_),
    .A2(_1643_),
    .B(_1089_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4723_ (.A1(_1245_),
    .A2(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4724_ (.A1(_1638_),
    .A2(_1721_),
    .B(_0948_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4725_ (.A1(_1717_),
    .A2(_1718_),
    .B(_3210_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4726_ (.A1(_1439_),
    .A2(_1268_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4727_ (.A1(_1277_),
    .A2(_1724_),
    .B(_0733_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4728_ (.A1(_1670_),
    .A2(_1558_),
    .B(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4729_ (.A1(_1072_),
    .A2(_1258_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4730_ (.A1(_1630_),
    .A2(_1727_),
    .B(_1073_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4731_ (.I0(_1309_),
    .I1(_1320_),
    .S(_1283_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4732_ (.A1(_1427_),
    .A2(_1542_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4733_ (.A1(_1670_),
    .A2(_1729_),
    .B(_1730_),
    .C(_1394_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4734_ (.A1(_1072_),
    .A2(_1501_),
    .B(_1728_),
    .C(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_1520_),
    .A2(_1726_),
    .B(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4736_ (.A1(_1719_),
    .A2(_1722_),
    .B(_1723_),
    .C(_1733_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4737_ (.A1(_1337_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4738_ (.A1(_1715_),
    .A2(_1735_),
    .B(_1518_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4739_ (.A1(_1351_),
    .A2(_1736_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4740_ (.A1(_0851_),
    .A2(_1336_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4741_ (.A1(_1347_),
    .A2(_1715_),
    .A3(_1735_),
    .B(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4742_ (.A1(_1518_),
    .A2(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4743_ (.A1(_1350_),
    .A2(_1737_),
    .B1(_1740_),
    .B2(_3212_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4744_ (.A1(_3194_),
    .A2(_3197_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4745_ (.I(_1742_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4746_ (.A1(_0727_),
    .A2(_1741_),
    .B(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4747_ (.I(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4748_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4749_ (.A1(_1346_),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4752_ (.I(_1050_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4753_ (.A1(_1750_),
    .A2(_1742_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4754_ (.I(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4755_ (.A1(\mod.pc_2[0] ),
    .A2(_1011_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4756_ (.A1(\mod.pc_2[0] ),
    .A2(_1011_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4757_ (.A1(_1752_),
    .A2(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4758_ (.A1(_1752_),
    .A2(_1344_),
    .B1(_1753_),
    .B2(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4759_ (.I(net13),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4760_ (.I(\mod.valid2 ),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4761_ (.I(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4762_ (.A1(_1750_),
    .A2(_3198_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4764_ (.A1(net15),
    .A2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4765_ (.A1(net14),
    .A2(_1760_),
    .B(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4766_ (.I(\mod.ldr_hzd[7] ),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4767_ (.I(\mod.ldr_hzd[6] ),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4768_ (.I(\mod.ldr_hzd[5] ),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4769_ (.I(\mod.ldr_hzd[4] ),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4770_ (.A1(_1764_),
    .A2(_1765_),
    .A3(_1766_),
    .A4(_1767_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(\mod.ldr_hzd[11] ),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4772_ (.I(\mod.ldr_hzd[10] ),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(\mod.ldr_hzd[9] ),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4774_ (.I(\mod.ldr_hzd[8] ),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4775_ (.A1(_1769_),
    .A2(_1770_),
    .A3(_1771_),
    .A4(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4776_ (.I(\mod.ldr_hzd[15] ),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4777_ (.I(\mod.ldr_hzd[14] ),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4778_ (.I(\mod.ldr_hzd[13] ),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4779_ (.I(\mod.ldr_hzd[12] ),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4780_ (.A1(_1774_),
    .A2(_1775_),
    .A3(_1776_),
    .A4(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(\mod.ldr_hzd[3] ),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4782_ (.I(\mod.ldr_hzd[2] ),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4783_ (.I(\mod.ldr_hzd[1] ),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4784_ (.I(\mod.ldr_hzd[0] ),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4785_ (.A1(_1779_),
    .A2(_1780_),
    .A3(_1781_),
    .A4(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4786_ (.A1(_1773_),
    .A2(_1778_),
    .A3(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4787_ (.I(_0977_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4788_ (.A1(_1765_),
    .A2(_1785_),
    .B(_0697_),
    .C(_0885_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_3133_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_0982_),
    .A2(_0445_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4791_ (.I(_3178_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4792_ (.A1(_1764_),
    .A2(_1787_),
    .B1(_1788_),
    .B2(_1766_),
    .C1(_1789_),
    .C2(_1767_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4793_ (.A1(_1786_),
    .A2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4794_ (.A1(_1774_),
    .A2(_1787_),
    .B(_0583_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4795_ (.A1(_1775_),
    .A2(_1785_),
    .B1(_1788_),
    .B2(_1776_),
    .C1(_1789_),
    .C2(_1777_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4796_ (.A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4797_ (.A1(_1782_),
    .A2(_1789_),
    .B(_0973_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4798_ (.A1(_1779_),
    .A2(_1787_),
    .B1(_1785_),
    .B2(_1780_),
    .C1(_1788_),
    .C2(_1781_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4799_ (.A1(_1772_),
    .A2(_1789_),
    .B(_0971_),
    .C(_0476_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4800_ (.A1(_1769_),
    .A2(_1787_),
    .B1(_1785_),
    .B2(_1770_),
    .C1(_1788_),
    .C2(_1771_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4801_ (.A1(_1795_),
    .A2(_1796_),
    .B1(_1797_),
    .B2(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4802_ (.A1(_1791_),
    .A2(_1794_),
    .A3(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4803_ (.I(_0609_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4804_ (.I(_0608_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4805_ (.I0(_1777_),
    .I1(_1776_),
    .I2(\mod.ldr_hzd[14] ),
    .I3(_1774_),
    .S0(_1801_),
    .S1(_1802_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4806_ (.A1(_0615_),
    .A2(_0607_),
    .A3(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4807_ (.I0(_1782_),
    .I1(\mod.ldr_hzd[1] ),
    .I2(\mod.ldr_hzd[2] ),
    .I3(\mod.ldr_hzd[3] ),
    .S0(_1801_),
    .S1(_1802_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4808_ (.A1(\mod.ldr_hzd[8] ),
    .A2(_0434_),
    .B(_0616_),
    .C(_0615_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4809_ (.A1(_1802_),
    .A2(_0429_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4810_ (.A1(_3236_),
    .A2(_1801_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4811_ (.A1(\mod.ldr_hzd[10] ),
    .A2(_1807_),
    .B1(_1808_),
    .B2(\mod.ldr_hzd[9] ),
    .C1(_0424_),
    .C2(\mod.ldr_hzd[11] ),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4812_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_1807_),
    .B(_0607_),
    .C(_0420_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4813_ (.A1(\mod.ldr_hzd[4] ),
    .A2(_0434_),
    .B1(_1808_),
    .B2(\mod.ldr_hzd[5] ),
    .C1(\mod.ldr_hzd[7] ),
    .C2(_0424_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4814_ (.A1(_1806_),
    .A2(_1809_),
    .B1(_1810_),
    .B2(_1811_),
    .C(_0944_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4815_ (.A1(_0613_),
    .A2(_1805_),
    .B(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4816_ (.A1(_1804_),
    .A2(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4817_ (.I(\mod.instr_2[6] ),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(\mod.instr_2[4] ),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4819_ (.I(\mod.instr_2[3] ),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4820_ (.I(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4821_ (.A1(_1816_),
    .A2(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_1819_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4823_ (.I(_1816_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4824_ (.A1(_1821_),
    .A2(_1818_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(_1822_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4826_ (.A1(_1781_),
    .A2(_1820_),
    .B1(_1823_),
    .B2(_1779_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4827_ (.A1(_1821_),
    .A2(_1817_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(_1825_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4829_ (.A1(_1816_),
    .A2(_1817_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4831_ (.A1(_1780_),
    .A2(_1826_),
    .B1(_1828_),
    .B2(\mod.ldr_hzd[0] ),
    .C(\mod.instr_2[5] ),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(_1824_),
    .A2(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(\mod.instr_2[5] ),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(_1765_),
    .A2(_1826_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4835_ (.A1(_1766_),
    .A2(_1820_),
    .B1(_1827_),
    .B2(_1767_),
    .C1(_1823_),
    .C2(_1764_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4836_ (.A1(_1831_),
    .A2(_1832_),
    .A3(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4837_ (.A1(_1815_),
    .A2(_1830_),
    .A3(_1834_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4838_ (.A1(_1775_),
    .A2(_1826_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4839_ (.A1(\mod.ldr_hzd[13] ),
    .A2(_1819_),
    .B1(_1827_),
    .B2(\mod.ldr_hzd[12] ),
    .C1(_1822_),
    .C2(\mod.ldr_hzd[15] ),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4840_ (.A1(_1831_),
    .A2(_1836_),
    .A3(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4841_ (.A1(_1771_),
    .A2(_1820_),
    .B1(_1823_),
    .B2(_1769_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4842_ (.A1(_1770_),
    .A2(_1825_),
    .B1(_1827_),
    .B2(_1772_),
    .C(\mod.instr_2[5] ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4843_ (.A1(_1839_),
    .A2(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4844_ (.A1(\mod.instr_2[6] ),
    .A2(_1838_),
    .A3(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4845_ (.A1(_1835_),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4846_ (.A1(_0729_),
    .A2(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4847_ (.A1(_0729_),
    .A2(_1800_),
    .B(_1814_),
    .C(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4848_ (.A1(_1768_),
    .A2(_1784_),
    .B(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4849_ (.A1(_1763_),
    .A2(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4850_ (.I(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4851_ (.A1(_1759_),
    .A2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4852_ (.I(\mod.valid0 ),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4853_ (.A1(_1745_),
    .A2(_1849_),
    .B(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4854_ (.A1(_1757_),
    .A2(_1851_),
    .B(_1848_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4856_ (.I(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4857_ (.A1(\mod.pc0[0] ),
    .A2(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4858_ (.I(net13),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4859_ (.A1(_0865_),
    .A2(_1349_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4860_ (.A1(_1351_),
    .A2(_1736_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4861_ (.A1(_0874_),
    .A2(_1739_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4862_ (.A1(_1857_),
    .A2(_1858_),
    .B1(_1859_),
    .B2(_1348_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4863_ (.A1(_3195_),
    .A2(_3196_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4864_ (.A1(_0728_),
    .A2(_1860_),
    .B(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4865_ (.A1(_1758_),
    .A2(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4866_ (.A1(_1850_),
    .A2(_1856_),
    .A3(_1863_),
    .B(_1847_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_1747_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_1866_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4870_ (.A1(\mod.pc[0] ),
    .A2(_1865_),
    .B(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4871_ (.A1(_1749_),
    .A2(_1756_),
    .B1(_1855_),
    .B2(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4872_ (.I(_3125_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4873_ (.A1(_3190_),
    .A2(_1344_),
    .B1(_1869_),
    .B2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(_3189_),
    .A2(_1871_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4875_ (.A1(\mod.des.des_counter[0] ),
    .A2(_3120_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4876_ (.I(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4877_ (.A1(_3211_),
    .A2(_1581_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4878_ (.I(_1864_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4879_ (.I(_1875_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4880_ (.A1(_1866_),
    .A2(_1875_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4881_ (.I(_1862_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4882_ (.I(\mod.pc[1] ),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4883_ (.A1(_1759_),
    .A2(_1878_),
    .B(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4884_ (.A1(\mod.pc0[1] ),
    .A2(_1876_),
    .B1(_1877_),
    .B2(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4885_ (.I(_1866_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4886_ (.I(_1861_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4887_ (.A1(_3200_),
    .A2(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_0992_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4889_ (.A1(_0830_),
    .A2(_1885_),
    .A3(_1753_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_1884_),
    .A2(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4891_ (.A1(_1884_),
    .A2(_1874_),
    .B(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4892_ (.A1(_1882_),
    .A2(_1888_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4893_ (.A1(_3126_),
    .A2(_1881_),
    .A3(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4894_ (.I(_3187_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4895_ (.A1(_0571_),
    .A2(_0592_),
    .B(_1891_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4896_ (.A1(_1873_),
    .A2(_1874_),
    .B(_1890_),
    .C(_1892_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_3210_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4898_ (.A1(_1893_),
    .A2(_1606_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4899_ (.I(_3125_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4900_ (.I(_1751_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4901_ (.I(\mod.pc_2[2] ),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4902_ (.I(_0961_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4903_ (.A1(_1038_),
    .A2(_1885_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_1038_),
    .A2(_1885_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4905_ (.A1(_1753_),
    .A2(_1899_),
    .B(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4906_ (.A1(_1897_),
    .A2(_1898_),
    .A3(_1901_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4907_ (.A1(_1896_),
    .A2(_1894_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4908_ (.A1(_1896_),
    .A2(_1902_),
    .B(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4909_ (.I(_1853_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4910_ (.A1(\mod.pc0[2] ),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4911_ (.A1(\mod.pc[2] ),
    .A2(_1865_),
    .B(_1867_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4912_ (.A1(_1749_),
    .A2(_1904_),
    .B1(_1906_),
    .B2(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4913_ (.A1(_1895_),
    .A2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_3188_),
    .A2(_1049_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4915_ (.A1(_1873_),
    .A2(_1894_),
    .B(_1909_),
    .C(_1910_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4916_ (.I(_1872_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4917_ (.A1(_1545_),
    .A2(_1564_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4918_ (.A1(_3211_),
    .A2(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4919_ (.I(_1105_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4920_ (.A1(_1897_),
    .A2(_1898_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4921_ (.A1(_1897_),
    .A2(_1898_),
    .B(_1901_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4922_ (.A1(_1915_),
    .A2(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4923_ (.A1(_1024_),
    .A2(_1914_),
    .A3(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4924_ (.A1(_1752_),
    .A2(_1913_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4925_ (.A1(_1896_),
    .A2(_1918_),
    .B(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4926_ (.A1(\mod.pc0[3] ),
    .A2(_1905_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4927_ (.A1(\mod.pc[3] ),
    .A2(_1865_),
    .B(_1748_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4928_ (.A1(_1749_),
    .A2(_1920_),
    .B1(_1921_),
    .B2(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4929_ (.A1(_1895_),
    .A2(_1923_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4930_ (.A1(_1891_),
    .A2(_1030_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4931_ (.A1(_1911_),
    .A2(_1913_),
    .B(_1924_),
    .C(_1925_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(_1884_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_1342_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4934_ (.A1(_1927_),
    .A2(_1538_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4935_ (.I(_1884_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4936_ (.A1(\mod.pc_2[4] ),
    .A2(_1122_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(\mod.pc_2[4] ),
    .A2(_1122_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4938_ (.A1(_1930_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4939_ (.A1(_1024_),
    .A2(_1914_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4940_ (.A1(_1024_),
    .A2(_1914_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4941_ (.A1(_1915_),
    .A2(_1933_),
    .A3(_1916_),
    .B(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4942_ (.A1(_1932_),
    .A2(_1935_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4943_ (.A1(_1929_),
    .A2(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4944_ (.A1(_1926_),
    .A2(_1928_),
    .B(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4945_ (.A1(\mod.pc0[4] ),
    .A2(_1854_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4946_ (.A1(\mod.pc[4] ),
    .A2(_1865_),
    .B(_1867_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4947_ (.A1(_1749_),
    .A2(_1938_),
    .B1(_1939_),
    .B2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4948_ (.A1(_1870_),
    .A2(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(_3190_),
    .A2(_1928_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4950_ (.A1(_0713_),
    .A2(_0719_),
    .B(_1891_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4951_ (.A1(_1942_),
    .A2(_1943_),
    .A3(_1944_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4952_ (.A1(_0000_),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4953_ (.A1(_1001_),
    .A2(_1002_),
    .A3(_1006_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4954_ (.I(_1758_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4955_ (.I(_1878_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4956_ (.A1(_1342_),
    .A2(_1522_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4957_ (.I(_1086_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4958_ (.I(_1931_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4959_ (.A1(_1930_),
    .A2(_1935_),
    .B(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4960_ (.A1(_0768_),
    .A2(_1950_),
    .A3(_1952_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4961_ (.A1(_1929_),
    .A2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4962_ (.A1(_1926_),
    .A2(_1949_),
    .B(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4963_ (.A1(_1947_),
    .A2(_1948_),
    .A3(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4964_ (.I(\mod.pc[5] ),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4965_ (.I(_1852_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4966_ (.A1(\mod.pc0[5] ),
    .A2(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_1863_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4968_ (.I(_1960_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4969_ (.A1(_1957_),
    .A2(_1854_),
    .B(_1959_),
    .C(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4970_ (.A1(_1956_),
    .A2(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4971_ (.A1(_3124_),
    .A2(_1949_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4972_ (.A1(_1945_),
    .A2(_1946_),
    .B1(_1963_),
    .B2(_0001_),
    .C(_1964_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4973_ (.I(_1759_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4974_ (.I(_1878_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4975_ (.A1(_1927_),
    .A2(_1635_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(\mod.pc_2[6] ),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4977_ (.I(_1070_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4978_ (.A1(_0768_),
    .A2(_1950_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4979_ (.A1(_1970_),
    .A2(_1952_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4980_ (.A1(_0768_),
    .A2(_1950_),
    .B(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4981_ (.A1(_1968_),
    .A2(_1969_),
    .A3(_1972_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4982_ (.A1(_1929_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4983_ (.A1(_1926_),
    .A2(_1967_),
    .B(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4984_ (.A1(_1965_),
    .A2(_1966_),
    .A3(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4985_ (.I(\mod.pc[6] ),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4986_ (.I(_1853_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4987_ (.A1(\mod.pc0[6] ),
    .A2(_1958_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4988_ (.I(_1960_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4989_ (.I(_1980_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4990_ (.A1(_1977_),
    .A2(_1978_),
    .B(_1979_),
    .C(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4991_ (.A1(_1976_),
    .A2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4992_ (.A1(_3124_),
    .A2(_1967_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_3187_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4994_ (.A1(_0970_),
    .A2(_0989_),
    .B(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4995_ (.A1(_3126_),
    .A2(_1983_),
    .B(_1984_),
    .C(_1986_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4996_ (.A1(_1700_),
    .A2(_1703_),
    .B(_1713_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4997_ (.A1(_3211_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4998_ (.I(_1752_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4999_ (.I(\mod.pc_2[7] ),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5000_ (.I(_0888_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5001_ (.I(_0890_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5002_ (.A1(_0586_),
    .A2(_1991_),
    .B(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5003_ (.A1(\mod.pc_2[6] ),
    .A2(_1969_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5004_ (.A1(_1968_),
    .A2(_1969_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5005_ (.A1(_1994_),
    .A2(_1972_),
    .B(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5006_ (.A1(_1990_),
    .A2(_1993_),
    .A3(_1996_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5007_ (.A1(_1896_),
    .A2(_1988_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5008_ (.A1(_1989_),
    .A2(_1997_),
    .B(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5009_ (.A1(_1947_),
    .A2(_1948_),
    .A3(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5010_ (.I(\mod.pc[7] ),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5011_ (.A1(\mod.pc0[7] ),
    .A2(_1853_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5012_ (.A1(_2001_),
    .A2(_1854_),
    .B(_2002_),
    .C(_1961_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5013_ (.A1(_2000_),
    .A2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5014_ (.A1(_0952_),
    .A2(_0957_),
    .B(_1985_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5015_ (.A1(_1911_),
    .A2(_1988_),
    .B1(_2004_),
    .B2(_0001_),
    .C(_2005_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5016_ (.A1(_1893_),
    .A2(_1485_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5017_ (.A1(_1098_),
    .A2(_1099_),
    .A3(_1103_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5018_ (.I(_1989_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5019_ (.A1(_0982_),
    .A2(_1991_),
    .B(_1992_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5020_ (.A1(_0663_),
    .A2(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5021_ (.A1(_0663_),
    .A2(_2009_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5022_ (.A1(_2010_),
    .A2(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5023_ (.A1(_1990_),
    .A2(_1993_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5024_ (.A1(_1990_),
    .A2(_1993_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5025_ (.A1(_2013_),
    .A2(_1996_),
    .B(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5026_ (.A1(_2012_),
    .A2(_2015_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5027_ (.A1(_1989_),
    .A2(_2006_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5028_ (.A1(_2008_),
    .A2(_2016_),
    .B(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5029_ (.A1(\mod.pc0[8] ),
    .A2(_1905_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5030_ (.A1(\mod.pc[8] ),
    .A2(_1875_),
    .B(_1748_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5031_ (.A1(_1882_),
    .A2(_2018_),
    .B1(_2019_),
    .B2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5032_ (.A1(_1891_),
    .A2(_2007_),
    .B1(_2021_),
    .B2(_1895_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5033_ (.A1(_1873_),
    .A2(_2006_),
    .B(_2022_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5034_ (.A1(_1927_),
    .A2(_1448_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5035_ (.I(\mod.pc_2[9] ),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5036_ (.A1(_0971_),
    .A2(_1991_),
    .B(_1992_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_2011_),
    .A2(_2015_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5038_ (.A1(_2010_),
    .A2(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5039_ (.A1(_2024_),
    .A2(_2025_),
    .A3(_2027_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5040_ (.A1(_1989_),
    .A2(_2023_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5041_ (.A1(_2008_),
    .A2(_2028_),
    .B(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5042_ (.A1(\mod.pc0[9] ),
    .A2(_1905_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5043_ (.A1(\mod.pc[9] ),
    .A2(_1875_),
    .B(_1748_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5044_ (.A1(_1882_),
    .A2(_2030_),
    .B1(_2031_),
    .B2(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5045_ (.A1(_1895_),
    .A2(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5046_ (.A1(_1115_),
    .A2(_1120_),
    .B(_1985_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5047_ (.A1(_1911_),
    .A2(_2023_),
    .B(_2034_),
    .C(_2035_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_1893_),
    .A2(_1659_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5049_ (.A1(\mod.pc0[10] ),
    .A2(_1958_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5050_ (.I(\mod.pc[10] ),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5051_ (.A1(_2038_),
    .A2(_1978_),
    .B(_1981_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5052_ (.I(_1929_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5053_ (.A1(_2024_),
    .A2(_2025_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5054_ (.A1(\mod.pc_2[9] ),
    .A2(_2025_),
    .B(_2027_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5055_ (.I(\mod.pc_2[10] ),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5056_ (.A1(_2043_),
    .A2(_0891_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5057_ (.A1(_2041_),
    .A2(_2042_),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5058_ (.A1(_2041_),
    .A2(_2044_),
    .A3(_2042_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_1926_),
    .A2(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5060_ (.A1(_2040_),
    .A2(_2036_),
    .B1(_2045_),
    .B2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5061_ (.A1(_1980_),
    .A2(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5062_ (.A1(_2037_),
    .A2(_2039_),
    .B(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5063_ (.A1(_1078_),
    .A2(_1083_),
    .B(_1985_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5064_ (.A1(_1911_),
    .A2(_2036_),
    .B1(_2050_),
    .B2(_0001_),
    .C(_2051_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5065_ (.I(_1927_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5066_ (.A1(_2052_),
    .A2(_1734_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_2008_),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5068_ (.A1(\mod.pc_2[10] ),
    .A2(_0891_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5069_ (.A1(_2055_),
    .A2(_2045_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5070_ (.I(\mod.pc_2[11] ),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5071_ (.I(\mod.funct7[0] ),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5072_ (.A1(_2058_),
    .A2(_1991_),
    .B(_1992_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5073_ (.A1(_2057_),
    .A2(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5074_ (.A1(_2056_),
    .A2(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5075_ (.A1(_2040_),
    .A2(_2061_),
    .B(_1966_),
    .C(_1965_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5076_ (.A1(\mod.pc0[11] ),
    .A2(_1958_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5077_ (.I(\mod.pc[11] ),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5078_ (.A1(_2064_),
    .A2(_1978_),
    .B(_1981_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5079_ (.A1(_2054_),
    .A2(_2062_),
    .B1(_2063_),
    .B2(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5080_ (.A1(_1064_),
    .A2(_1068_),
    .B(_3187_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5081_ (.A1(_1872_),
    .A2(_2053_),
    .B1(_2066_),
    .B2(_3126_),
    .C(_2067_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5082_ (.A1(_2052_),
    .A2(_1406_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5083_ (.A1(\mod.pc_2[12] ),
    .A2(_1177_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5084_ (.A1(_2057_),
    .A2(_2059_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5085_ (.A1(_2055_),
    .A2(_2045_),
    .B(_2060_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5086_ (.A1(_2070_),
    .A2(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5087_ (.A1(_2069_),
    .A2(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5088_ (.I0(_2068_),
    .I1(_2073_),
    .S(_2040_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5089_ (.A1(_1981_),
    .A2(_2074_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5090_ (.I(\mod.pc0[12] ),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5091_ (.A1(\mod.pc[12] ),
    .A2(_1866_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5092_ (.A1(_2076_),
    .A2(_1876_),
    .B1(_1877_),
    .B2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5093_ (.A1(_2075_),
    .A2(_2078_),
    .B(_1870_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5094_ (.A1(_3188_),
    .A2(_1152_),
    .B1(_2068_),
    .B2(_3190_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5095_ (.A1(_2079_),
    .A2(_2080_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5096_ (.A1(_1893_),
    .A2(_1679_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(_3190_),
    .A2(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5098_ (.A1(\mod.pc0[13] ),
    .A2(_1978_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5099_ (.A1(\mod.pc[13] ),
    .A2(_1876_),
    .B(_1867_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5100_ (.I(_1177_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_2069_),
    .A2(_2072_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5102_ (.A1(_1138_),
    .A2(_2085_),
    .B(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5103_ (.A1(_1209_),
    .A2(_2085_),
    .A3(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5104_ (.A1(_2040_),
    .A2(_2081_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5105_ (.A1(_2008_),
    .A2(_2088_),
    .B(_2089_),
    .C(_1961_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5106_ (.A1(_2083_),
    .A2(_2084_),
    .B(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5107_ (.A1(_3188_),
    .A2(_1168_),
    .B1(_2091_),
    .B2(_1870_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(_2082_),
    .A2(_2092_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5109_ (.A1(_2052_),
    .A2(_1694_),
    .A3(_1697_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5110_ (.A1(_1945_),
    .A2(_1190_),
    .B1(_2093_),
    .B2(_1873_),
    .ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5111_ (.A1(_1760_),
    .A2(_1849_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_2094_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5113_ (.A1(_1347_),
    .A2(net22),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5114_ (.I(_2095_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5115_ (.I(net11),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_2096_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5117_ (.I(_2097_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5118_ (.I(_1831_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5119_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5120_ (.I(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5121_ (.I(_2099_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5122_ (.A1(\mod.rd_3[2] ),
    .A2(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5123_ (.A1(_2098_),
    .A2(_2100_),
    .B(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5124_ (.I(_1815_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5125_ (.I(_2099_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(\mod.rd_3[3] ),
    .A2(_2100_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5127_ (.A1(_2104_),
    .A2(_2105_),
    .B(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5128_ (.A1(_2103_),
    .A2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5129_ (.I(net12),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5130_ (.A1(_2109_),
    .A2(_1848_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5131_ (.A1(\mod.valid2 ),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5132_ (.A1(net12),
    .A2(_2101_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5133_ (.A1(_0944_),
    .A2(_2111_),
    .B(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5134_ (.I(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5135_ (.A1(\mod.rd_3[1] ),
    .A2(_2101_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5136_ (.A1(_1821_),
    .A2(_2100_),
    .B(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(\mod.rd_3[0] ),
    .A2(_2101_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5138_ (.A1(_1818_),
    .A2(_2100_),
    .B(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5139_ (.I(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5140_ (.A1(_2114_),
    .A2(_2116_),
    .A3(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_2108_),
    .A2(_2120_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5142_ (.I(_2121_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5143_ (.I(_2122_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5144_ (.I(_2105_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5145_ (.I(_2124_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5146_ (.I(_1883_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5147_ (.I(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5148_ (.A1(_2126_),
    .A2(_1344_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5149_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5150_ (.A1(_1750_),
    .A2(_3201_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(_2129_),
    .A2(_2130_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5152_ (.I(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5153_ (.A1(_3224_),
    .A2(_2127_),
    .B(_2128_),
    .C(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5154_ (.A1(\mod.des.des_dout[21] ),
    .A2(_2125_),
    .B(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5155_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5156_ (.I(_2121_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5157_ (.I(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5158_ (.A1(\mod.registers.r1[0] ),
    .A2(_2137_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5159_ (.A1(_2123_),
    .A2(_2135_),
    .B(_2138_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5160_ (.I(_1743_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5161_ (.I(_1743_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5162_ (.A1(_1038_),
    .A2(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5163_ (.A1(_2139_),
    .A2(_1874_),
    .B(_2132_),
    .C(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5164_ (.A1(\mod.des.des_dout[22] ),
    .A2(_2125_),
    .B(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5165_ (.I(_2143_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5166_ (.A1(\mod.registers.r1[1] ),
    .A2(_2137_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5167_ (.A1(_2123_),
    .A2(_2144_),
    .B(_2145_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5168_ (.A1(_1897_),
    .A2(_2140_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5169_ (.A1(_2139_),
    .A2(_1894_),
    .B(_2132_),
    .C(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5170_ (.A1(\mod.des.des_dout[23] ),
    .A2(_2125_),
    .B(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5171_ (.I(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5172_ (.A1(\mod.registers.r1[2] ),
    .A2(_2137_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5173_ (.A1(_2123_),
    .A2(_2149_),
    .B(_2150_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5174_ (.I(_2124_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5175_ (.I(_1743_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5176_ (.A1(_2152_),
    .A2(_1913_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5177_ (.I(_2126_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5178_ (.I(_2131_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5179_ (.A1(_0799_),
    .A2(_2154_),
    .B(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5180_ (.A1(\mod.des.des_dout[24] ),
    .A2(_2151_),
    .B1(_2153_),
    .B2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5181_ (.I(_2157_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5182_ (.A1(\mod.registers.r1[3] ),
    .A2(_2137_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5183_ (.A1(_2123_),
    .A2(_2158_),
    .B(_2159_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5184_ (.I(_2122_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(\mod.pc_2[4] ),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5186_ (.A1(_2126_),
    .A2(_1928_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5187_ (.A1(_2161_),
    .A2(_2127_),
    .B(_2132_),
    .C(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5188_ (.A1(\mod.des.des_dout[25] ),
    .A2(_2125_),
    .B(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5189_ (.I(_2164_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5190_ (.I(_2136_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(\mod.registers.r1[4] ),
    .A2(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5192_ (.A1(_2160_),
    .A2(_2165_),
    .B(_2167_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5193_ (.I(_2130_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5194_ (.A1(_2139_),
    .A2(_1949_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5195_ (.A1(_0769_),
    .A2(_2152_),
    .B(_2168_),
    .C(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5196_ (.I(_2105_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5197_ (.I(_2130_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5198_ (.A1(_1011_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5199_ (.A1(_2171_),
    .A2(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5200_ (.A1(\mod.des.des_dout[26] ),
    .A2(_2151_),
    .B1(_2170_),
    .B2(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5201_ (.I(_2175_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(\mod.registers.r1[5] ),
    .A2(_2166_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5203_ (.A1(_2160_),
    .A2(_2176_),
    .B(_2177_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5204_ (.I(_2129_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5205_ (.I(_1883_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5206_ (.A1(_2179_),
    .A2(_1967_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5207_ (.I(_2130_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5208_ (.A1(_1968_),
    .A2(_2139_),
    .B(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5209_ (.A1(_3200_),
    .A2(_0934_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5210_ (.A1(_1885_),
    .A2(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5211_ (.I(_2129_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5212_ (.A1(_2180_),
    .A2(_2182_),
    .B(_2184_),
    .C(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5213_ (.A1(\mod.des.des_dout[27] ),
    .A2(_2178_),
    .B(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5214_ (.I(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5215_ (.A1(\mod.registers.r1[6] ),
    .A2(_2166_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5216_ (.A1(_2160_),
    .A2(_2188_),
    .B(_2189_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5217_ (.A1(_1990_),
    .A2(_2179_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5218_ (.A1(_2154_),
    .A2(_1988_),
    .B(_2168_),
    .C(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5219_ (.A1(_1898_),
    .A2(_2172_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5220_ (.A1(_2171_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5221_ (.A1(\mod.des.des_dout[28] ),
    .A2(_2151_),
    .B1(_2191_),
    .B2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5222_ (.I(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5223_ (.A1(\mod.registers.r1[7] ),
    .A2(_2166_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5224_ (.A1(_2160_),
    .A2(_2195_),
    .B(_2196_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5225_ (.I(_2122_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5226_ (.I(_1883_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5227_ (.A1(_0663_),
    .A2(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5228_ (.A1(_2154_),
    .A2(_2006_),
    .B(_2168_),
    .C(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5229_ (.A1(_1914_),
    .A2(_2172_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5230_ (.A1(_2171_),
    .A2(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5231_ (.A1(\mod.des.des_dout[29] ),
    .A2(_2151_),
    .B1(_2200_),
    .B2(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5232_ (.I(_2203_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5233_ (.I(_2136_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(\mod.registers.r1[8] ),
    .A2(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5235_ (.A1(_2197_),
    .A2(_2204_),
    .B(_2206_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5236_ (.I(_2105_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5237_ (.I(_2181_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(_2024_),
    .A2(_2198_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5239_ (.A1(_2154_),
    .A2(_2023_),
    .B(_2208_),
    .C(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5240_ (.A1(_1122_),
    .A2(_2181_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5241_ (.A1(_2124_),
    .A2(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5242_ (.A1(\mod.des.des_dout[30] ),
    .A2(_2207_),
    .B1(_2210_),
    .B2(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5243_ (.I(_2213_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(\mod.registers.r1[9] ),
    .A2(_2205_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5245_ (.A1(_2197_),
    .A2(_2214_),
    .B(_2215_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5246_ (.A1(\mod.pc_2[10] ),
    .A2(_2198_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5247_ (.A1(_2127_),
    .A2(_2036_),
    .B(_2208_),
    .C(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5248_ (.A1(_1950_),
    .A2(_2185_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(_2155_),
    .A2(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5250_ (.A1(\mod.des.des_dout[31] ),
    .A2(_2207_),
    .B1(_2217_),
    .B2(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_2220_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(\mod.registers.r1[10] ),
    .A2(_2205_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5253_ (.A1(_2197_),
    .A2(_2221_),
    .B(_2222_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(_2057_),
    .A2(_2198_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5255_ (.A1(_2127_),
    .A2(_2053_),
    .B(_2208_),
    .C(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5256_ (.A1(_1969_),
    .A2(_2181_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5257_ (.A1(_2124_),
    .A2(_2225_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5258_ (.A1(\mod.des.des_dout[32] ),
    .A2(_2207_),
    .B1(_2224_),
    .B2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5259_ (.I(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5260_ (.A1(\mod.registers.r1[11] ),
    .A2(_2205_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5261_ (.A1(_2197_),
    .A2(_2228_),
    .B(_2229_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5262_ (.I(_2122_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5263_ (.A1(_2140_),
    .A2(_2068_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5264_ (.A1(_1138_),
    .A2(_2152_),
    .B(_2208_),
    .C(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5265_ (.A1(_1993_),
    .A2(_2185_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(_2155_),
    .A2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5267_ (.A1(\mod.des.des_dout[33] ),
    .A2(_2207_),
    .B1(_2232_),
    .B2(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5268_ (.I(_2235_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5269_ (.I(_2136_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5270_ (.A1(\mod.registers.r1[12] ),
    .A2(_2237_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5271_ (.A1(_2230_),
    .A2(_2236_),
    .B(_2238_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5272_ (.A1(_2140_),
    .A2(_2081_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5273_ (.A1(_1209_),
    .A2(_2152_),
    .B(_2172_),
    .C(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_2009_),
    .A2(_2129_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(_2155_),
    .A2(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5276_ (.A1(\mod.des.des_dout[34] ),
    .A2(_2171_),
    .B1(_2240_),
    .B2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5277_ (.I(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(\mod.registers.r1[13] ),
    .A2(_2237_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5279_ (.A1(_2230_),
    .A2(_2244_),
    .B(_2245_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5280_ (.A1(_2179_),
    .A2(_2093_),
    .A3(_2183_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5281_ (.A1(_1179_),
    .A2(_2168_),
    .B(_2185_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5282_ (.A1(\mod.des.des_dout[35] ),
    .A2(_2178_),
    .B1(_2246_),
    .B2(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5283_ (.I(_2248_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(\mod.registers.r1[14] ),
    .A2(_2237_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5285_ (.A1(_2230_),
    .A2(_2249_),
    .B(_2250_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5286_ (.A1(_2179_),
    .A2(_2052_),
    .A3(_1337_),
    .A4(_2183_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5287_ (.A1(_0891_),
    .A2(_2183_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5288_ (.A1(_2178_),
    .A2(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5289_ (.A1(\mod.des.des_dout[36] ),
    .A2(_2178_),
    .B1(_2251_),
    .B2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5290_ (.I(_2254_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5291_ (.A1(\mod.registers.r1[15] ),
    .A2(_2237_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5292_ (.A1(_2230_),
    .A2(_2255_),
    .B(_2256_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(_2113_),
    .A2(_2116_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5294_ (.A1(_2118_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5295_ (.A1(_2108_),
    .A2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5296_ (.I(_2259_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5297_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5298_ (.I(_2259_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5299_ (.I(_2262_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5300_ (.A1(\mod.registers.r2[0] ),
    .A2(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5301_ (.A1(_2135_),
    .A2(_2261_),
    .B(_2264_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(\mod.registers.r2[1] ),
    .A2(_2263_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5303_ (.A1(_2144_),
    .A2(_2261_),
    .B(_2265_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5304_ (.A1(\mod.registers.r2[2] ),
    .A2(_2263_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5305_ (.A1(_2149_),
    .A2(_2261_),
    .B(_2266_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5306_ (.A1(\mod.registers.r2[3] ),
    .A2(_2263_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5307_ (.A1(_2158_),
    .A2(_2261_),
    .B(_2267_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5308_ (.I(_2260_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5309_ (.I(_2262_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(\mod.registers.r2[4] ),
    .A2(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5311_ (.A1(_2165_),
    .A2(_2268_),
    .B(_2270_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5312_ (.A1(\mod.registers.r2[5] ),
    .A2(_2269_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5313_ (.A1(_2176_),
    .A2(_2268_),
    .B(_2271_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5314_ (.A1(\mod.registers.r2[6] ),
    .A2(_2269_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5315_ (.A1(_2188_),
    .A2(_2268_),
    .B(_2272_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5316_ (.A1(\mod.registers.r2[7] ),
    .A2(_2269_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5317_ (.A1(_2195_),
    .A2(_2268_),
    .B(_2273_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5318_ (.I(_2260_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5319_ (.I(_2262_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5320_ (.A1(\mod.registers.r2[8] ),
    .A2(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5321_ (.A1(_2204_),
    .A2(_2274_),
    .B(_2276_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5322_ (.A1(\mod.registers.r2[9] ),
    .A2(_2275_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(_2214_),
    .A2(_2274_),
    .B(_2277_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5324_ (.A1(\mod.registers.r2[10] ),
    .A2(_2275_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5325_ (.A1(_2221_),
    .A2(_2274_),
    .B(_2278_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5326_ (.A1(\mod.registers.r2[11] ),
    .A2(_2275_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5327_ (.A1(_2228_),
    .A2(_2274_),
    .B(_2279_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_2260_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_2262_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5330_ (.A1(\mod.registers.r2[12] ),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5331_ (.A1(_2236_),
    .A2(_2280_),
    .B(_2282_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(\mod.registers.r2[13] ),
    .A2(_2281_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5333_ (.A1(_2244_),
    .A2(_2280_),
    .B(_2283_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5334_ (.A1(\mod.registers.r2[14] ),
    .A2(_2281_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5335_ (.A1(_2249_),
    .A2(_2280_),
    .B(_2284_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(\mod.registers.r2[15] ),
    .A2(_2281_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5337_ (.A1(_2255_),
    .A2(_2280_),
    .B(_2285_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5338_ (.A1(_2119_),
    .A2(_2257_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5339_ (.A1(_2108_),
    .A2(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5340_ (.I(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5341_ (.I(_2288_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_2287_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_2290_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5344_ (.A1(\mod.registers.r3[0] ),
    .A2(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5345_ (.A1(_2135_),
    .A2(_2289_),
    .B(_2292_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5346_ (.A1(\mod.registers.r3[1] ),
    .A2(_2291_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5347_ (.A1(_2144_),
    .A2(_2289_),
    .B(_2293_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5348_ (.A1(\mod.registers.r3[2] ),
    .A2(_2291_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5349_ (.A1(_2149_),
    .A2(_2289_),
    .B(_2294_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5350_ (.A1(\mod.registers.r3[3] ),
    .A2(_2291_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5351_ (.A1(_2158_),
    .A2(_2289_),
    .B(_2295_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5352_ (.I(_2288_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_2290_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5354_ (.A1(\mod.registers.r3[4] ),
    .A2(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5355_ (.A1(_2165_),
    .A2(_2296_),
    .B(_2298_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5356_ (.A1(\mod.registers.r3[5] ),
    .A2(_2297_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5357_ (.A1(_2176_),
    .A2(_2296_),
    .B(_2299_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5358_ (.A1(\mod.registers.r3[6] ),
    .A2(_2297_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5359_ (.A1(_2188_),
    .A2(_2296_),
    .B(_2300_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5360_ (.A1(\mod.registers.r3[7] ),
    .A2(_2297_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5361_ (.A1(_2195_),
    .A2(_2296_),
    .B(_2301_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(_2288_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5363_ (.I(_2290_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5364_ (.A1(\mod.registers.r3[8] ),
    .A2(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5365_ (.A1(_2204_),
    .A2(_2302_),
    .B(_2304_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5366_ (.A1(\mod.registers.r3[9] ),
    .A2(_2303_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5367_ (.A1(_2214_),
    .A2(_2302_),
    .B(_2305_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5368_ (.A1(\mod.registers.r3[10] ),
    .A2(_2303_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5369_ (.A1(_2221_),
    .A2(_2302_),
    .B(_2306_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5370_ (.A1(\mod.registers.r3[11] ),
    .A2(_2303_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5371_ (.A1(_2228_),
    .A2(_2302_),
    .B(_2307_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5372_ (.I(_2288_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_2290_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5374_ (.A1(\mod.registers.r3[12] ),
    .A2(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5375_ (.A1(_2236_),
    .A2(_2308_),
    .B(_2310_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5376_ (.A1(\mod.registers.r3[13] ),
    .A2(_2309_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5377_ (.A1(_2244_),
    .A2(_2308_),
    .B(_2311_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5378_ (.A1(\mod.registers.r3[14] ),
    .A2(_2309_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5379_ (.A1(_2249_),
    .A2(_2308_),
    .B(_2312_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(\mod.registers.r3[15] ),
    .A2(_2309_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5381_ (.A1(_2255_),
    .A2(_2308_),
    .B(_2313_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5382_ (.I(_2103_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5383_ (.A1(_2314_),
    .A2(_2107_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5384_ (.A1(_2114_),
    .A2(_2116_),
    .A3(_2118_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5385_ (.A1(_2315_),
    .A2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5386_ (.I(_2317_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5387_ (.I(_2318_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5388_ (.I(_2317_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5389_ (.I(_2320_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5390_ (.A1(\mod.registers.r4[0] ),
    .A2(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5391_ (.A1(_2135_),
    .A2(_2319_),
    .B(_2322_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(\mod.registers.r4[1] ),
    .A2(_2321_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5393_ (.A1(_2144_),
    .A2(_2319_),
    .B(_2323_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5394_ (.A1(\mod.registers.r4[2] ),
    .A2(_2321_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5395_ (.A1(_2149_),
    .A2(_2319_),
    .B(_2324_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5396_ (.A1(\mod.registers.r4[3] ),
    .A2(_2321_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5397_ (.A1(_2158_),
    .A2(_2319_),
    .B(_2325_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5398_ (.I(_2318_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5399_ (.I(_2320_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5400_ (.A1(\mod.registers.r4[4] ),
    .A2(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5401_ (.A1(_2165_),
    .A2(_2326_),
    .B(_2328_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(\mod.registers.r4[5] ),
    .A2(_2327_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5403_ (.A1(_2176_),
    .A2(_2326_),
    .B(_2329_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(\mod.registers.r4[6] ),
    .A2(_2327_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5405_ (.A1(_2188_),
    .A2(_2326_),
    .B(_2330_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5406_ (.A1(\mod.registers.r4[7] ),
    .A2(_2327_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5407_ (.A1(_2195_),
    .A2(_2326_),
    .B(_2331_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(_2318_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_2320_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5410_ (.A1(\mod.registers.r4[8] ),
    .A2(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5411_ (.A1(_2204_),
    .A2(_2332_),
    .B(_2334_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5412_ (.A1(\mod.registers.r4[9] ),
    .A2(_2333_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5413_ (.A1(_2214_),
    .A2(_2332_),
    .B(_2335_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(\mod.registers.r4[10] ),
    .A2(_2333_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5415_ (.A1(_2221_),
    .A2(_2332_),
    .B(_2336_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(\mod.registers.r4[11] ),
    .A2(_2333_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5417_ (.A1(_2228_),
    .A2(_2332_),
    .B(_2337_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5418_ (.I(_2318_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5419_ (.I(_2320_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(\mod.registers.r4[12] ),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(_2236_),
    .A2(_2338_),
    .B(_2340_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5422_ (.A1(\mod.registers.r4[13] ),
    .A2(_2339_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5423_ (.A1(_2244_),
    .A2(_2338_),
    .B(_2341_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(\mod.registers.r4[14] ),
    .A2(_2339_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5425_ (.A1(_2249_),
    .A2(_2338_),
    .B(_2342_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5426_ (.A1(\mod.registers.r4[15] ),
    .A2(_2339_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5427_ (.A1(_2255_),
    .A2(_2338_),
    .B(_2343_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_2134_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5429_ (.I(_2344_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(_2120_),
    .A2(_2315_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5431_ (.I(_2346_),
    .Z(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_2347_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5433_ (.I(_2346_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5434_ (.I(_2349_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5435_ (.A1(\mod.registers.r5[0] ),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5436_ (.A1(_2345_),
    .A2(_2348_),
    .B(_2351_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5437_ (.I(_2143_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5438_ (.I(_2352_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5439_ (.A1(\mod.registers.r5[1] ),
    .A2(_2350_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5440_ (.A1(_2353_),
    .A2(_2348_),
    .B(_2354_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_2148_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5442_ (.I(_2355_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5443_ (.A1(\mod.registers.r5[2] ),
    .A2(_2350_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5444_ (.A1(_2356_),
    .A2(_2348_),
    .B(_2357_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5445_ (.I(_2157_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5446_ (.I(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5447_ (.A1(\mod.registers.r5[3] ),
    .A2(_2350_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5448_ (.A1(_2359_),
    .A2(_2348_),
    .B(_2360_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5449_ (.I(_2164_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5450_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5451_ (.I(_2347_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5452_ (.I(_2349_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(\mod.registers.r5[4] ),
    .A2(_2364_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5454_ (.A1(_2362_),
    .A2(_2363_),
    .B(_2365_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5455_ (.I(_2175_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5456_ (.I(_2366_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5457_ (.A1(\mod.registers.r5[5] ),
    .A2(_2364_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5458_ (.A1(_2367_),
    .A2(_2363_),
    .B(_2368_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_2187_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5460_ (.I(_2369_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5461_ (.A1(\mod.registers.r5[6] ),
    .A2(_2364_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5462_ (.A1(_2370_),
    .A2(_2363_),
    .B(_2371_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5463_ (.I(_2194_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5464_ (.I(_2372_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5465_ (.A1(\mod.registers.r5[7] ),
    .A2(_2364_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5466_ (.A1(_2373_),
    .A2(_2363_),
    .B(_2374_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5467_ (.I(_2203_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5468_ (.I(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_2347_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_2349_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5471_ (.A1(\mod.registers.r5[8] ),
    .A2(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5472_ (.A1(_2376_),
    .A2(_2377_),
    .B(_2379_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5473_ (.I(_2213_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5474_ (.I(_2380_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5475_ (.A1(\mod.registers.r5[9] ),
    .A2(_2378_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5476_ (.A1(_2381_),
    .A2(_2377_),
    .B(_2382_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5477_ (.I(_2220_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5478_ (.I(_2383_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5479_ (.A1(\mod.registers.r5[10] ),
    .A2(_2378_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5480_ (.A1(_2384_),
    .A2(_2377_),
    .B(_2385_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5481_ (.I(_2227_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5482_ (.I(_2386_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5483_ (.A1(\mod.registers.r5[11] ),
    .A2(_2378_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5484_ (.A1(_2387_),
    .A2(_2377_),
    .B(_2388_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5485_ (.I(_2235_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5486_ (.I(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5487_ (.I(_2347_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5488_ (.I(_2349_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(\mod.registers.r5[12] ),
    .A2(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5490_ (.A1(_2390_),
    .A2(_2391_),
    .B(_2393_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5491_ (.I(_2243_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5492_ (.I(_2394_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5493_ (.A1(\mod.registers.r5[13] ),
    .A2(_2392_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5494_ (.A1(_2395_),
    .A2(_2391_),
    .B(_2396_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5495_ (.I(_2248_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5496_ (.I(_2397_),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5497_ (.A1(\mod.registers.r5[14] ),
    .A2(_2392_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5498_ (.A1(_2398_),
    .A2(_2391_),
    .B(_2399_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_2254_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5500_ (.I(_2400_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5501_ (.A1(\mod.registers.r5[15] ),
    .A2(_2392_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5502_ (.A1(_2401_),
    .A2(_2391_),
    .B(_2402_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5503_ (.A1(_2258_),
    .A2(_2315_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5504_ (.I(_2403_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5505_ (.I(_2404_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5506_ (.I(_2403_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5507_ (.I(_2406_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5508_ (.A1(\mod.registers.r6[0] ),
    .A2(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5509_ (.A1(_2345_),
    .A2(_2405_),
    .B(_2408_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(\mod.registers.r6[1] ),
    .A2(_2407_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5511_ (.A1(_2353_),
    .A2(_2405_),
    .B(_2409_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(\mod.registers.r6[2] ),
    .A2(_2407_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5513_ (.A1(_2356_),
    .A2(_2405_),
    .B(_2410_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5514_ (.A1(\mod.registers.r6[3] ),
    .A2(_2407_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5515_ (.A1(_2359_),
    .A2(_2405_),
    .B(_2411_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5516_ (.I(_2404_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5517_ (.I(_2406_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5518_ (.A1(\mod.registers.r6[4] ),
    .A2(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5519_ (.A1(_2362_),
    .A2(_2412_),
    .B(_2414_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(\mod.registers.r6[5] ),
    .A2(_2413_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_2367_),
    .A2(_2412_),
    .B(_2415_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5522_ (.A1(\mod.registers.r6[6] ),
    .A2(_2413_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5523_ (.A1(_2370_),
    .A2(_2412_),
    .B(_2416_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5524_ (.A1(\mod.registers.r6[7] ),
    .A2(_2413_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5525_ (.A1(_2373_),
    .A2(_2412_),
    .B(_2417_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5526_ (.I(_2404_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5527_ (.I(_2406_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5528_ (.A1(\mod.registers.r6[8] ),
    .A2(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5529_ (.A1(_2376_),
    .A2(_2418_),
    .B(_2420_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5530_ (.A1(\mod.registers.r6[9] ),
    .A2(_2419_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5531_ (.A1(_2381_),
    .A2(_2418_),
    .B(_2421_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5532_ (.A1(\mod.registers.r6[10] ),
    .A2(_2419_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5533_ (.A1(_2384_),
    .A2(_2418_),
    .B(_2422_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(\mod.registers.r6[11] ),
    .A2(_2419_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5535_ (.A1(_2387_),
    .A2(_2418_),
    .B(_2423_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5536_ (.I(_2404_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5537_ (.I(_2406_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5538_ (.A1(\mod.registers.r6[12] ),
    .A2(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5539_ (.A1(_2390_),
    .A2(_2424_),
    .B(_2426_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5540_ (.A1(\mod.registers.r6[13] ),
    .A2(_2425_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5541_ (.A1(_2395_),
    .A2(_2424_),
    .B(_2427_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5542_ (.A1(\mod.registers.r6[14] ),
    .A2(_2425_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5543_ (.A1(_2398_),
    .A2(_2424_),
    .B(_2428_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5544_ (.A1(\mod.registers.r6[15] ),
    .A2(_2425_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5545_ (.A1(_2401_),
    .A2(_2424_),
    .B(_2429_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5546_ (.A1(_2286_),
    .A2(_2315_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5547_ (.I(_2430_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5548_ (.I(_2431_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5549_ (.I(_2430_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5550_ (.I(_2433_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(\mod.registers.r7[0] ),
    .A2(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5552_ (.A1(_2345_),
    .A2(_2432_),
    .B(_2435_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5553_ (.A1(\mod.registers.r7[1] ),
    .A2(_2434_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5554_ (.A1(_2353_),
    .A2(_2432_),
    .B(_2436_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5555_ (.A1(\mod.registers.r7[2] ),
    .A2(_2434_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5556_ (.A1(_2356_),
    .A2(_2432_),
    .B(_2437_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5557_ (.A1(\mod.registers.r7[3] ),
    .A2(_2434_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5558_ (.A1(_2359_),
    .A2(_2432_),
    .B(_2438_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5559_ (.I(_2431_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5560_ (.I(_2433_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5561_ (.A1(\mod.registers.r7[4] ),
    .A2(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5562_ (.A1(_2362_),
    .A2(_2439_),
    .B(_2441_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5563_ (.A1(\mod.registers.r7[5] ),
    .A2(_2440_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5564_ (.A1(_2367_),
    .A2(_2439_),
    .B(_2442_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5565_ (.A1(\mod.registers.r7[6] ),
    .A2(_2440_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5566_ (.A1(_2370_),
    .A2(_2439_),
    .B(_2443_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5567_ (.A1(\mod.registers.r7[7] ),
    .A2(_2440_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5568_ (.A1(_2373_),
    .A2(_2439_),
    .B(_2444_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_2431_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5570_ (.I(_2433_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5571_ (.A1(\mod.registers.r7[8] ),
    .A2(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5572_ (.A1(_2376_),
    .A2(_2445_),
    .B(_2447_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5573_ (.A1(\mod.registers.r7[9] ),
    .A2(_2446_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5574_ (.A1(_2381_),
    .A2(_2445_),
    .B(_2448_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5575_ (.A1(\mod.registers.r7[10] ),
    .A2(_2446_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5576_ (.A1(_2384_),
    .A2(_2445_),
    .B(_2449_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5577_ (.A1(\mod.registers.r7[11] ),
    .A2(_2446_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5578_ (.A1(_2387_),
    .A2(_2445_),
    .B(_2450_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_2431_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5580_ (.I(_2433_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5581_ (.A1(\mod.registers.r7[12] ),
    .A2(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5582_ (.A1(_2390_),
    .A2(_2451_),
    .B(_2453_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5583_ (.A1(\mod.registers.r7[13] ),
    .A2(_2452_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5584_ (.A1(_2395_),
    .A2(_2451_),
    .B(_2454_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5585_ (.A1(\mod.registers.r7[14] ),
    .A2(_2452_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5586_ (.A1(_2398_),
    .A2(_2451_),
    .B(_2455_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5587_ (.A1(\mod.registers.r7[15] ),
    .A2(_2452_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5588_ (.A1(_2401_),
    .A2(_2451_),
    .B(_2456_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5589_ (.I(_2107_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5590_ (.A1(_2103_),
    .A2(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5591_ (.A1(_2316_),
    .A2(_2458_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_2459_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5593_ (.I(_2460_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5594_ (.I(_2459_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5595_ (.I(_2462_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5596_ (.A1(\mod.registers.r8[0] ),
    .A2(_2463_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5597_ (.A1(_2345_),
    .A2(_2461_),
    .B(_2464_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(\mod.registers.r8[1] ),
    .A2(_2463_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5599_ (.A1(_2353_),
    .A2(_2461_),
    .B(_2465_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5600_ (.A1(\mod.registers.r8[2] ),
    .A2(_2463_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5601_ (.A1(_2356_),
    .A2(_2461_),
    .B(_2466_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5602_ (.A1(\mod.registers.r8[3] ),
    .A2(_2463_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5603_ (.A1(_2359_),
    .A2(_2461_),
    .B(_2467_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5604_ (.I(_2460_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5605_ (.I(_2462_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5606_ (.A1(\mod.registers.r8[4] ),
    .A2(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5607_ (.A1(_2362_),
    .A2(_2468_),
    .B(_2470_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5608_ (.A1(\mod.registers.r8[5] ),
    .A2(_2469_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5609_ (.A1(_2367_),
    .A2(_2468_),
    .B(_2471_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5610_ (.A1(\mod.registers.r8[6] ),
    .A2(_2469_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5611_ (.A1(_2370_),
    .A2(_2468_),
    .B(_2472_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5612_ (.A1(\mod.registers.r8[7] ),
    .A2(_2469_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5613_ (.A1(_2373_),
    .A2(_2468_),
    .B(_2473_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_2460_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5615_ (.I(_2462_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5616_ (.A1(\mod.registers.r8[8] ),
    .A2(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5617_ (.A1(_2376_),
    .A2(_2474_),
    .B(_2476_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5618_ (.A1(\mod.registers.r8[9] ),
    .A2(_2475_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5619_ (.A1(_2381_),
    .A2(_2474_),
    .B(_2477_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5620_ (.A1(\mod.registers.r8[10] ),
    .A2(_2475_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5621_ (.A1(_2384_),
    .A2(_2474_),
    .B(_2478_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5622_ (.A1(\mod.registers.r8[11] ),
    .A2(_2475_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5623_ (.A1(_2387_),
    .A2(_2474_),
    .B(_2479_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5624_ (.I(_2460_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(_2462_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5626_ (.A1(\mod.registers.r8[12] ),
    .A2(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5627_ (.A1(_2390_),
    .A2(_2480_),
    .B(_2482_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5628_ (.A1(\mod.registers.r8[13] ),
    .A2(_2481_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5629_ (.A1(_2395_),
    .A2(_2480_),
    .B(_2483_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(\mod.registers.r8[14] ),
    .A2(_2481_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5631_ (.A1(_2398_),
    .A2(_2480_),
    .B(_2484_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5632_ (.A1(\mod.registers.r8[15] ),
    .A2(_2481_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5633_ (.A1(_2401_),
    .A2(_2480_),
    .B(_2485_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5634_ (.I(_2134_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5635_ (.A1(_2120_),
    .A2(_2458_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5636_ (.I(_2487_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5638_ (.I(_2487_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5639_ (.I(_2490_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5640_ (.A1(\mod.registers.r9[0] ),
    .A2(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5641_ (.A1(_2486_),
    .A2(_2489_),
    .B(_2492_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5642_ (.I(_2143_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5643_ (.A1(\mod.registers.r9[1] ),
    .A2(_2491_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_2493_),
    .A2(_2489_),
    .B(_2494_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5645_ (.I(_2148_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5646_ (.A1(\mod.registers.r9[2] ),
    .A2(_2491_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5647_ (.A1(_2495_),
    .A2(_2489_),
    .B(_2496_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5648_ (.I(_2157_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5649_ (.A1(\mod.registers.r9[3] ),
    .A2(_2491_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5650_ (.A1(_2497_),
    .A2(_2489_),
    .B(_2498_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5651_ (.I(_2164_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5652_ (.I(_2488_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_2490_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5654_ (.A1(\mod.registers.r9[4] ),
    .A2(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5655_ (.A1(_2499_),
    .A2(_2500_),
    .B(_2502_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5656_ (.I(_2175_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\mod.registers.r9[5] ),
    .A2(_2501_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_2503_),
    .A2(_2500_),
    .B(_2504_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_2187_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5660_ (.A1(\mod.registers.r9[6] ),
    .A2(_2501_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5661_ (.A1(_2505_),
    .A2(_2500_),
    .B(_2506_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5662_ (.I(_2194_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(\mod.registers.r9[7] ),
    .A2(_2501_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5664_ (.A1(_2507_),
    .A2(_2500_),
    .B(_2508_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_2203_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5666_ (.I(_2488_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5667_ (.I(_2490_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(\mod.registers.r9[8] ),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5669_ (.A1(_2509_),
    .A2(_2510_),
    .B(_2512_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5670_ (.I(_2213_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5671_ (.A1(\mod.registers.r9[9] ),
    .A2(_2511_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5672_ (.A1(_2513_),
    .A2(_2510_),
    .B(_2514_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(_2220_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5674_ (.A1(\mod.registers.r9[10] ),
    .A2(_2511_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_2515_),
    .A2(_2510_),
    .B(_2516_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5676_ (.I(_2227_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5677_ (.A1(\mod.registers.r9[11] ),
    .A2(_2511_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5678_ (.A1(_2517_),
    .A2(_2510_),
    .B(_2518_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5679_ (.I(_2235_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5680_ (.I(_2488_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5681_ (.I(_2490_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5682_ (.A1(\mod.registers.r9[12] ),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5683_ (.A1(_2519_),
    .A2(_2520_),
    .B(_2522_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5684_ (.I(_2243_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5685_ (.A1(\mod.registers.r9[13] ),
    .A2(_2521_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5686_ (.A1(_2523_),
    .A2(_2520_),
    .B(_2524_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_2248_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(\mod.registers.r9[14] ),
    .A2(_2521_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(_2525_),
    .A2(_2520_),
    .B(_2526_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_2254_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5691_ (.A1(\mod.registers.r9[15] ),
    .A2(_2521_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5692_ (.A1(_2527_),
    .A2(_2520_),
    .B(_2528_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5693_ (.A1(_2258_),
    .A2(_2458_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_2529_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_2530_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5696_ (.I(_2529_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5697_ (.I(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5698_ (.A1(\mod.registers.r10[0] ),
    .A2(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_2486_),
    .A2(_2531_),
    .B(_2534_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5700_ (.A1(\mod.registers.r10[1] ),
    .A2(_2533_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5701_ (.A1(_2493_),
    .A2(_2531_),
    .B(_2535_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5702_ (.A1(\mod.registers.r10[2] ),
    .A2(_2533_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5703_ (.A1(_2495_),
    .A2(_2531_),
    .B(_2536_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5704_ (.A1(\mod.registers.r10[3] ),
    .A2(_2533_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5705_ (.A1(_2497_),
    .A2(_2531_),
    .B(_2537_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_2530_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_2532_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5708_ (.A1(\mod.registers.r10[4] ),
    .A2(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5709_ (.A1(_2499_),
    .A2(_2538_),
    .B(_2540_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(\mod.registers.r10[5] ),
    .A2(_2539_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5711_ (.A1(_2503_),
    .A2(_2538_),
    .B(_2541_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(\mod.registers.r10[6] ),
    .A2(_2539_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5713_ (.A1(_2505_),
    .A2(_2538_),
    .B(_2542_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5714_ (.A1(\mod.registers.r10[7] ),
    .A2(_2539_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5715_ (.A1(_2507_),
    .A2(_2538_),
    .B(_2543_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5716_ (.I(_2530_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5717_ (.I(_2532_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(\mod.registers.r10[8] ),
    .A2(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5719_ (.A1(_2509_),
    .A2(_2544_),
    .B(_2546_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5720_ (.A1(\mod.registers.r10[9] ),
    .A2(_2545_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5721_ (.A1(_2513_),
    .A2(_2544_),
    .B(_2547_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5722_ (.A1(\mod.registers.r10[10] ),
    .A2(_2545_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5723_ (.A1(_2515_),
    .A2(_2544_),
    .B(_2548_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5724_ (.A1(\mod.registers.r10[11] ),
    .A2(_2545_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5725_ (.A1(_2517_),
    .A2(_2544_),
    .B(_2549_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5726_ (.I(_2530_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_2532_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5728_ (.A1(\mod.registers.r10[12] ),
    .A2(_2551_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5729_ (.A1(_2519_),
    .A2(_2550_),
    .B(_2552_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(\mod.registers.r10[13] ),
    .A2(_2551_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5731_ (.A1(_2523_),
    .A2(_2550_),
    .B(_2553_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5732_ (.A1(\mod.registers.r10[14] ),
    .A2(_2551_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5733_ (.A1(_2525_),
    .A2(_2550_),
    .B(_2554_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5734_ (.A1(\mod.registers.r10[15] ),
    .A2(_2551_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5735_ (.A1(_2527_),
    .A2(_2550_),
    .B(_2555_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5736_ (.A1(_2286_),
    .A2(_2458_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_2556_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5738_ (.I(_2557_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5739_ (.I(_2556_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5740_ (.I(_2559_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5741_ (.A1(\mod.registers.r11[0] ),
    .A2(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5742_ (.A1(_2486_),
    .A2(_2558_),
    .B(_2561_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5743_ (.A1(\mod.registers.r11[1] ),
    .A2(_2560_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5744_ (.A1(_2493_),
    .A2(_2558_),
    .B(_2562_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(\mod.registers.r11[2] ),
    .A2(_2560_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5746_ (.A1(_2495_),
    .A2(_2558_),
    .B(_2563_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5747_ (.A1(\mod.registers.r11[3] ),
    .A2(_2560_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5748_ (.A1(_2497_),
    .A2(_2558_),
    .B(_2564_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_2557_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(_2559_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5751_ (.A1(\mod.registers.r11[4] ),
    .A2(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5752_ (.A1(_2499_),
    .A2(_2565_),
    .B(_2567_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(\mod.registers.r11[5] ),
    .A2(_2566_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5754_ (.A1(_2503_),
    .A2(_2565_),
    .B(_2568_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5755_ (.A1(\mod.registers.r11[6] ),
    .A2(_2566_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5756_ (.A1(_2505_),
    .A2(_2565_),
    .B(_2569_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5757_ (.A1(\mod.registers.r11[7] ),
    .A2(_2566_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5758_ (.A1(_2507_),
    .A2(_2565_),
    .B(_2570_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5759_ (.I(_2557_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_2559_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5761_ (.A1(\mod.registers.r11[8] ),
    .A2(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5762_ (.A1(_2509_),
    .A2(_2571_),
    .B(_2573_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5763_ (.A1(\mod.registers.r11[9] ),
    .A2(_2572_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5764_ (.A1(_2513_),
    .A2(_2571_),
    .B(_2574_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5765_ (.A1(\mod.registers.r11[10] ),
    .A2(_2572_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5766_ (.A1(_2515_),
    .A2(_2571_),
    .B(_2575_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5767_ (.A1(\mod.registers.r11[11] ),
    .A2(_2572_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5768_ (.A1(_2517_),
    .A2(_2571_),
    .B(_2576_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5769_ (.I(_2557_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5770_ (.I(_2559_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5771_ (.A1(\mod.registers.r11[12] ),
    .A2(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5772_ (.A1(_2519_),
    .A2(_2577_),
    .B(_2579_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5773_ (.A1(\mod.registers.r11[13] ),
    .A2(_2578_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5774_ (.A1(_2523_),
    .A2(_2577_),
    .B(_2580_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5775_ (.A1(\mod.registers.r11[14] ),
    .A2(_2578_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5776_ (.A1(_2525_),
    .A2(_2577_),
    .B(_2581_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5777_ (.A1(\mod.registers.r11[15] ),
    .A2(_2578_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5778_ (.A1(_2527_),
    .A2(_2577_),
    .B(_2582_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5779_ (.A1(_2314_),
    .A2(_2457_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5780_ (.A1(_2316_),
    .A2(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5781_ (.I(_2584_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5782_ (.I(_2585_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5783_ (.I(_2584_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5784_ (.I(_2587_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(\mod.registers.r12[0] ),
    .A2(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5786_ (.A1(_2486_),
    .A2(_2586_),
    .B(_2589_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(\mod.registers.r12[1] ),
    .A2(_2588_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5788_ (.A1(_2493_),
    .A2(_2586_),
    .B(_2590_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5789_ (.A1(\mod.registers.r12[2] ),
    .A2(_2588_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5790_ (.A1(_2495_),
    .A2(_2586_),
    .B(_2591_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5791_ (.A1(\mod.registers.r12[3] ),
    .A2(_2588_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5792_ (.A1(_2497_),
    .A2(_2586_),
    .B(_2592_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_2585_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5794_ (.I(_2587_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5795_ (.A1(\mod.registers.r12[4] ),
    .A2(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5796_ (.A1(_2499_),
    .A2(_2593_),
    .B(_2595_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(\mod.registers.r12[5] ),
    .A2(_2594_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5798_ (.A1(_2503_),
    .A2(_2593_),
    .B(_2596_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5799_ (.A1(\mod.registers.r12[6] ),
    .A2(_2594_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5800_ (.A1(_2505_),
    .A2(_2593_),
    .B(_2597_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5801_ (.A1(\mod.registers.r12[7] ),
    .A2(_2594_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5802_ (.A1(_2507_),
    .A2(_2593_),
    .B(_2598_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(_2585_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5804_ (.I(_2587_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5805_ (.A1(\mod.registers.r12[8] ),
    .A2(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5806_ (.A1(_2509_),
    .A2(_2599_),
    .B(_2601_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(\mod.registers.r12[9] ),
    .A2(_2600_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5808_ (.A1(_2513_),
    .A2(_2599_),
    .B(_2602_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5809_ (.A1(\mod.registers.r12[10] ),
    .A2(_2600_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5810_ (.A1(_2515_),
    .A2(_2599_),
    .B(_2603_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(\mod.registers.r12[11] ),
    .A2(_2600_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5812_ (.A1(_2517_),
    .A2(_2599_),
    .B(_2604_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5813_ (.I(_2585_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5814_ (.I(_2587_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(\mod.registers.r12[12] ),
    .A2(_2606_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5816_ (.A1(_2519_),
    .A2(_2605_),
    .B(_2607_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(\mod.registers.r12[13] ),
    .A2(_2606_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(_2523_),
    .A2(_2605_),
    .B(_2608_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5819_ (.A1(\mod.registers.r12[14] ),
    .A2(_2606_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5820_ (.A1(_2525_),
    .A2(_2605_),
    .B(_2609_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5821_ (.A1(\mod.registers.r12[15] ),
    .A2(_2606_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5822_ (.A1(_2527_),
    .A2(_2605_),
    .B(_2610_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5823_ (.A1(_2120_),
    .A2(_2583_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5824_ (.I(_2611_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5825_ (.I(_2612_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5826_ (.I(_2611_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5827_ (.I(_2614_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(\mod.registers.r13[0] ),
    .A2(_2615_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5829_ (.A1(_2344_),
    .A2(_2613_),
    .B(_2616_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5830_ (.A1(\mod.registers.r13[1] ),
    .A2(_2615_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5831_ (.A1(_2352_),
    .A2(_2613_),
    .B(_2617_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5832_ (.A1(\mod.registers.r13[2] ),
    .A2(_2615_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5833_ (.A1(_2355_),
    .A2(_2613_),
    .B(_2618_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(\mod.registers.r13[3] ),
    .A2(_2615_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5835_ (.A1(_2358_),
    .A2(_2613_),
    .B(_2619_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5836_ (.I(_2612_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5837_ (.I(_2614_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5838_ (.A1(\mod.registers.r13[4] ),
    .A2(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5839_ (.A1(_2361_),
    .A2(_2620_),
    .B(_2622_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(\mod.registers.r13[5] ),
    .A2(_2621_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5841_ (.A1(_2366_),
    .A2(_2620_),
    .B(_2623_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(\mod.registers.r13[6] ),
    .A2(_2621_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5843_ (.A1(_2369_),
    .A2(_2620_),
    .B(_2624_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5844_ (.A1(\mod.registers.r13[7] ),
    .A2(_2621_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5845_ (.A1(_2372_),
    .A2(_2620_),
    .B(_2625_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5846_ (.I(_2612_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5847_ (.I(_2614_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5848_ (.A1(\mod.registers.r13[8] ),
    .A2(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5849_ (.A1(_2375_),
    .A2(_2626_),
    .B(_2628_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5850_ (.A1(\mod.registers.r13[9] ),
    .A2(_2627_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5851_ (.A1(_2380_),
    .A2(_2626_),
    .B(_2629_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5852_ (.A1(\mod.registers.r13[10] ),
    .A2(_2627_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5853_ (.A1(_2383_),
    .A2(_2626_),
    .B(_2630_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5854_ (.A1(\mod.registers.r13[11] ),
    .A2(_2627_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5855_ (.A1(_2386_),
    .A2(_2626_),
    .B(_2631_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5856_ (.I(_2612_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5857_ (.I(_2614_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5858_ (.A1(\mod.registers.r13[12] ),
    .A2(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5859_ (.A1(_2389_),
    .A2(_2632_),
    .B(_2634_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5860_ (.A1(\mod.registers.r13[13] ),
    .A2(_2633_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5861_ (.A1(_2394_),
    .A2(_2632_),
    .B(_2635_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5862_ (.A1(\mod.registers.r13[14] ),
    .A2(_2633_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5863_ (.A1(_2397_),
    .A2(_2632_),
    .B(_2636_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5864_ (.A1(\mod.registers.r13[15] ),
    .A2(_2633_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5865_ (.A1(_2400_),
    .A2(_2632_),
    .B(_2637_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5866_ (.A1(_2258_),
    .A2(_2583_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5867_ (.I(_2638_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5868_ (.I(_2639_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5869_ (.I(_2638_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_2641_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5871_ (.A1(\mod.registers.r14[0] ),
    .A2(_2642_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5872_ (.A1(_2344_),
    .A2(_2640_),
    .B(_2643_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5873_ (.A1(\mod.registers.r14[1] ),
    .A2(_2642_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5874_ (.A1(_2352_),
    .A2(_2640_),
    .B(_2644_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5875_ (.A1(\mod.registers.r14[2] ),
    .A2(_2642_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5876_ (.A1(_2355_),
    .A2(_2640_),
    .B(_2645_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5877_ (.A1(\mod.registers.r14[3] ),
    .A2(_2642_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5878_ (.A1(_2358_),
    .A2(_2640_),
    .B(_2646_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5879_ (.I(_2639_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5880_ (.I(_2641_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5881_ (.A1(\mod.registers.r14[4] ),
    .A2(_2648_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5882_ (.A1(_2361_),
    .A2(_2647_),
    .B(_2649_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5883_ (.A1(\mod.registers.r14[5] ),
    .A2(_2648_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5884_ (.A1(_2366_),
    .A2(_2647_),
    .B(_2650_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5885_ (.A1(\mod.registers.r14[6] ),
    .A2(_2648_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5886_ (.A1(_2369_),
    .A2(_2647_),
    .B(_2651_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5887_ (.A1(\mod.registers.r14[7] ),
    .A2(_2648_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5888_ (.A1(_2372_),
    .A2(_2647_),
    .B(_2652_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_2639_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5890_ (.I(_2641_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(\mod.registers.r14[8] ),
    .A2(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5892_ (.A1(_2375_),
    .A2(_2653_),
    .B(_2655_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(\mod.registers.r14[9] ),
    .A2(_2654_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5894_ (.A1(_2380_),
    .A2(_2653_),
    .B(_2656_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(\mod.registers.r14[10] ),
    .A2(_2654_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5896_ (.A1(_2383_),
    .A2(_2653_),
    .B(_2657_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(\mod.registers.r14[11] ),
    .A2(_2654_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5898_ (.A1(_2386_),
    .A2(_2653_),
    .B(_2658_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5899_ (.I(_2639_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5900_ (.I(_2641_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5901_ (.A1(\mod.registers.r14[12] ),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5902_ (.A1(_2389_),
    .A2(_2659_),
    .B(_2661_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5903_ (.A1(\mod.registers.r14[13] ),
    .A2(_2660_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5904_ (.A1(_2394_),
    .A2(_2659_),
    .B(_2662_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5905_ (.A1(\mod.registers.r14[14] ),
    .A2(_2660_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5906_ (.A1(_2397_),
    .A2(_2659_),
    .B(_2663_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5907_ (.A1(\mod.registers.r14[15] ),
    .A2(_2660_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5908_ (.A1(_2400_),
    .A2(_2659_),
    .B(_2664_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5909_ (.I(net11),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5910_ (.I(_2665_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_2666_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5912_ (.I(_2667_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5913_ (.I(_2667_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5914_ (.I(_2667_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5915_ (.I(_2110_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5916_ (.I(_2668_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5917_ (.I(_2669_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_1851_),
    .A2(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5920_ (.A1(_2667_),
    .A2(_2672_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5921_ (.A1(_1851_),
    .A2(_2668_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5922_ (.I(_2673_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5923_ (.I(_2674_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5924_ (.I(net12),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5925_ (.A1(_2676_),
    .A2(_1847_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5926_ (.I(_2677_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_2678_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5928_ (.I(\mod.valid1 ),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5929_ (.A1(_1746_),
    .A2(_1849_),
    .B(_2680_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(_2679_),
    .A2(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5931_ (.I(_2665_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5932_ (.I(_2683_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5933_ (.A1(_2675_),
    .A2(_2682_),
    .B(_2684_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5934_ (.I(_2676_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5935_ (.A1(_2685_),
    .A2(\mod.pc0[0] ),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5936_ (.I(_2109_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5937_ (.I(_2687_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5938_ (.A1(_2688_),
    .A2(_1869_),
    .B(_0003_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5939_ (.A1(_2686_),
    .A2(_2689_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_2676_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5941_ (.A1(_1881_),
    .A2(_1889_),
    .B(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5942_ (.A1(_2690_),
    .A2(\mod.pc0[1] ),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5943_ (.A1(_0003_),
    .A2(_2691_),
    .A3(_2692_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5944_ (.I(_2693_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5945_ (.A1(_2685_),
    .A2(\mod.pc0[2] ),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5946_ (.I(_2096_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(_2695_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5948_ (.A1(_2688_),
    .A2(_1908_),
    .B(_2696_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5949_ (.A1(_2694_),
    .A2(_2697_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_2676_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5951_ (.I(_2698_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5952_ (.A1(_2699_),
    .A2(\mod.pc0[3] ),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5953_ (.A1(_2688_),
    .A2(_1923_),
    .B(_2696_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5954_ (.A1(_2700_),
    .A2(_2701_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5955_ (.A1(_2699_),
    .A2(\mod.pc0[4] ),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5956_ (.I(_2687_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5957_ (.A1(_2703_),
    .A2(_1941_),
    .B(_2696_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5958_ (.A1(_2702_),
    .A2(_2704_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_2690_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_2698_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5961_ (.I(_2695_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5962_ (.A1(_2706_),
    .A2(\mod.pc0[5] ),
    .B(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5963_ (.A1(_2705_),
    .A2(_1963_),
    .B(_2708_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5964_ (.A1(_2706_),
    .A2(\mod.pc0[6] ),
    .B(_2707_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5965_ (.A1(_2705_),
    .A2(_1983_),
    .B(_2709_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5966_ (.I(_2695_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5967_ (.A1(_2706_),
    .A2(\mod.pc0[7] ),
    .B(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5968_ (.A1(_2705_),
    .A2(_2004_),
    .B(_2711_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5969_ (.A1(_2699_),
    .A2(\mod.pc0[8] ),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5970_ (.A1(_2703_),
    .A2(_2021_),
    .B(_2696_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5971_ (.A1(_2712_),
    .A2(_2713_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5972_ (.A1(_2699_),
    .A2(\mod.pc0[9] ),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5973_ (.A1(_2703_),
    .A2(_2033_),
    .B(_2707_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5974_ (.A1(_2714_),
    .A2(_2715_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5975_ (.A1(_2706_),
    .A2(\mod.pc0[10] ),
    .B(_2710_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5976_ (.A1(_2705_),
    .A2(_2050_),
    .B(_2716_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5977_ (.A1(_2690_),
    .A2(\mod.pc0[11] ),
    .B(_2710_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5978_ (.A1(_2685_),
    .A2(_2066_),
    .B(_2717_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(net11),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5980_ (.I(_2718_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5981_ (.A1(_2687_),
    .A2(_2075_),
    .A3(_2078_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5982_ (.A1(_2688_),
    .A2(_2076_),
    .B(_2719_),
    .C(_2720_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5983_ (.A1(\mod.pc0[13] ),
    .A2(_2685_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5984_ (.A1(_2703_),
    .A2(_2091_),
    .B(_2707_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5985_ (.A1(_2721_),
    .A2(_2722_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5986_ (.A1(_1747_),
    .A2(_1864_),
    .B(_2109_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5987_ (.I(_2723_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5988_ (.I(_2724_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5989_ (.A1(_1947_),
    .A2(_1948_),
    .A3(_1756_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5990_ (.I(\mod.pc[0] ),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5991_ (.A1(_1345_),
    .A2(_1745_),
    .B(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5992_ (.A1(_2726_),
    .A2(_2728_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5993_ (.I(_2723_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5994_ (.A1(\mod.pc[0] ),
    .A2(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5995_ (.I(_2718_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5996_ (.A1(_2725_),
    .A2(_2729_),
    .B(_2731_),
    .C(_2732_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5997_ (.I(_2730_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5998_ (.A1(_1759_),
    .A2(_1878_),
    .A3(_1888_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5999_ (.A1(_1880_),
    .A2(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6000_ (.A1(_2729_),
    .A2(_2735_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_2724_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6002_ (.A1(\mod.pc[1] ),
    .A2(_2737_),
    .B(_2710_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6003_ (.A1(_2733_),
    .A2(_2736_),
    .B(_2738_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6004_ (.A1(_2726_),
    .A2(_2728_),
    .B(_1880_),
    .C(_2734_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6005_ (.I(_2739_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6006_ (.A1(_1965_),
    .A2(_1966_),
    .A3(_1904_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6007_ (.I(\mod.valid2 ),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6008_ (.I(_1744_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6009_ (.I(\mod.pc[2] ),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6010_ (.A1(_2742_),
    .A2(_2743_),
    .B(_2744_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6011_ (.A1(_2741_),
    .A2(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6012_ (.A1(_2740_),
    .A2(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6013_ (.I(_2695_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6014_ (.A1(\mod.pc[2] ),
    .A2(_2737_),
    .B(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6015_ (.A1(_2733_),
    .A2(_2747_),
    .B(_2749_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6016_ (.I(\mod.pc[3] ),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6017_ (.A1(_2698_),
    .A2(_1877_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6018_ (.I(_2751_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6019_ (.A1(_1947_),
    .A2(_1948_),
    .A3(_1920_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6020_ (.A1(_1345_),
    .A2(_2743_),
    .B(_2750_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6021_ (.A1(_2741_),
    .A2(_2745_),
    .B1(_2753_),
    .B2(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6022_ (.A1(_2740_),
    .A2(_2755_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6023_ (.I(_2756_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6024_ (.A1(_2753_),
    .A2(_2754_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6025_ (.A1(_2740_),
    .A2(_2746_),
    .B(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6026_ (.A1(_2757_),
    .A2(_2759_),
    .B(_2751_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6027_ (.A1(_2750_),
    .A2(_2752_),
    .B(_2760_),
    .C(_2719_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6028_ (.A1(_1965_),
    .A2(_1966_),
    .A3(_1938_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6029_ (.I(\mod.pc[4] ),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6030_ (.A1(_2742_),
    .A2(_2743_),
    .B(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6031_ (.A1(_2761_),
    .A2(_2763_),
    .Z(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6032_ (.A1(_2757_),
    .A2(_2764_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6033_ (.I(_2723_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6034_ (.A1(\mod.pc[4] ),
    .A2(_2766_),
    .B(_2748_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6035_ (.A1(_2733_),
    .A2(_2765_),
    .B(_2767_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6036_ (.A1(_2740_),
    .A2(_2755_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6037_ (.A1(_1345_),
    .A2(_1745_),
    .B(_1957_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6038_ (.A1(_2768_),
    .A2(_2764_),
    .B(_1956_),
    .C(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6039_ (.A1(_2761_),
    .A2(_2763_),
    .B1(_1956_),
    .B2(_2769_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6040_ (.A1(_2756_),
    .A2(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6041_ (.A1(_2770_),
    .A2(_2772_),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6042_ (.A1(\mod.pc[5] ),
    .A2(_2724_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6043_ (.A1(_2737_),
    .A2(_2773_),
    .B(_2774_),
    .C(_2719_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6044_ (.A1(_2742_),
    .A2(_1746_),
    .B(_1977_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6045_ (.A1(_1976_),
    .A2(_2775_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6046_ (.A1(_2772_),
    .A2(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6047_ (.A1(\mod.pc[6] ),
    .A2(_2766_),
    .B(_2748_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6048_ (.A1(_2733_),
    .A2(_2777_),
    .B(_2778_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6049_ (.A1(\mod.pc[7] ),
    .A2(_2752_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6050_ (.A1(_2742_),
    .A2(_2743_),
    .B(_2001_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6051_ (.A1(_2757_),
    .A2(_2771_),
    .A3(_2776_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6052_ (.A1(_1976_),
    .A2(_2775_),
    .B1(_2000_),
    .B2(_2780_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6053_ (.A1(_2739_),
    .A2(_2755_),
    .A3(_2771_),
    .A4(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6054_ (.I(_2783_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6055_ (.A1(_1882_),
    .A2(_1876_),
    .B(_2784_),
    .C(_2687_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6056_ (.A1(_2000_),
    .A2(_2780_),
    .A3(_2781_),
    .B(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6057_ (.A1(_2779_),
    .A2(_2786_),
    .B(_2684_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6058_ (.I(\mod.pc[8] ),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6059_ (.I0(_2787_),
    .I1(_2018_),
    .S(_1960_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6060_ (.A1(_2784_),
    .A2(_2788_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6061_ (.A1(\mod.pc[8] ),
    .A2(_2766_),
    .B(_2748_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6062_ (.A1(_2725_),
    .A2(_2789_),
    .B(_2790_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6063_ (.A1(\mod.pc[9] ),
    .A2(_2752_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6064_ (.A1(_2757_),
    .A2(_2771_),
    .A3(_2782_),
    .A4(_2788_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6065_ (.I(\mod.pc[9] ),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6066_ (.I0(_2793_),
    .I1(_2030_),
    .S(_1960_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6067_ (.I(_2794_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6068_ (.A1(_2788_),
    .A2(_2794_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6069_ (.A1(_2783_),
    .A2(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6070_ (.A1(_2792_),
    .A2(_2795_),
    .B(_2797_),
    .C(_2730_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6071_ (.I(_2666_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6072_ (.A1(_2791_),
    .A2(_2798_),
    .B(_2799_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6073_ (.A1(_1346_),
    .A2(_1746_),
    .B(_2038_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6074_ (.A1(_2049_),
    .A2(_2800_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6075_ (.A1(_2797_),
    .A2(_2801_),
    .Z(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6076_ (.A1(\mod.pc[10] ),
    .A2(_2724_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6077_ (.A1(_2737_),
    .A2(_2802_),
    .B(_2803_),
    .C(_2719_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6078_ (.A1(_2784_),
    .A2(_2796_),
    .A3(_2801_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6079_ (.A1(\mod.pc[11] ),
    .A2(_1747_),
    .B1(_2054_),
    .B2(_2062_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6080_ (.I(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6081_ (.A1(_1980_),
    .A2(_2048_),
    .B(_2800_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6082_ (.A1(_2788_),
    .A2(_2794_),
    .A3(_2807_),
    .A4(_2805_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6083_ (.A1(_2783_),
    .A2(_2808_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6084_ (.A1(_2804_),
    .A2(_2806_),
    .B(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6085_ (.I(_2096_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6086_ (.I(_2811_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6087_ (.A1(\mod.pc[11] ),
    .A2(_2766_),
    .B(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6088_ (.A1(_2725_),
    .A2(_2810_),
    .B(_2813_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6089_ (.A1(_1980_),
    .A2(_2074_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6090_ (.A1(_2814_),
    .A2(_2077_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6091_ (.A1(_2809_),
    .A2(_2815_),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6092_ (.A1(\mod.pc[12] ),
    .A2(_2730_),
    .B(_2812_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6093_ (.A1(_2725_),
    .A2(_2816_),
    .B(_2817_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6094_ (.I(\mod.pc[13] ),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6095_ (.A1(_2784_),
    .A2(_2808_),
    .A3(_2815_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6096_ (.A1(_2818_),
    .A2(_1961_),
    .B(_2090_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6097_ (.A1(_2819_),
    .A2(_2820_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6098_ (.A1(_2819_),
    .A2(_2820_),
    .B(_2751_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(_2683_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6100_ (.A1(_2818_),
    .A2(_2752_),
    .B1(_2821_),
    .B2(_2822_),
    .C(_2823_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_2669_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6102_ (.I(_2824_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6103_ (.I(_2669_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6104_ (.I(_2826_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6105_ (.A1(\mod.pc_1[0] ),
    .A2(_2827_),
    .B(_2812_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6106_ (.A1(_2727_),
    .A2(_2825_),
    .B(_2828_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6107_ (.A1(\mod.pc_1[1] ),
    .A2(_2827_),
    .B(_2812_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6108_ (.A1(_1879_),
    .A2(_2825_),
    .B(_2829_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_2811_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6110_ (.A1(\mod.pc_1[2] ),
    .A2(_2827_),
    .B(_2830_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6111_ (.A1(_2744_),
    .A2(_2825_),
    .B(_2831_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6112_ (.A1(\mod.pc_1[3] ),
    .A2(_2827_),
    .B(_2830_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6113_ (.A1(_2750_),
    .A2(_2825_),
    .B(_2832_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6114_ (.I(_2824_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6115_ (.I(_2826_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6116_ (.A1(\mod.pc_1[4] ),
    .A2(_2834_),
    .B(_2830_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6117_ (.A1(_2762_),
    .A2(_2833_),
    .B(_2835_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6118_ (.A1(\mod.pc_1[5] ),
    .A2(_2834_),
    .B(_2830_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6119_ (.A1(_1957_),
    .A2(_2833_),
    .B(_2836_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6120_ (.I(_2811_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6121_ (.A1(\mod.pc_1[6] ),
    .A2(_2834_),
    .B(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6122_ (.A1(_1977_),
    .A2(_2833_),
    .B(_2838_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6123_ (.A1(\mod.pc_1[7] ),
    .A2(_2834_),
    .B(_2837_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6124_ (.A1(_2001_),
    .A2(_2833_),
    .B(_2839_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6125_ (.I(_2670_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6126_ (.I(_2826_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6127_ (.A1(\mod.pc_1[8] ),
    .A2(_2841_),
    .B(_2837_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6128_ (.A1(_2787_),
    .A2(_2840_),
    .B(_2842_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6129_ (.A1(\mod.pc_1[9] ),
    .A2(_2841_),
    .B(_2837_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6130_ (.A1(_2793_),
    .A2(_2840_),
    .B(_2843_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6131_ (.I(_2811_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6132_ (.A1(\mod.pc_1[10] ),
    .A2(_2841_),
    .B(_2844_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6133_ (.A1(_2038_),
    .A2(_2840_),
    .B(_2845_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6134_ (.A1(\mod.pc_1[11] ),
    .A2(_2841_),
    .B(_2844_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6135_ (.A1(_2064_),
    .A2(_2840_),
    .B(_2846_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6136_ (.I(\mod.pc_1[12] ),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6137_ (.I(_2677_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6138_ (.I(_2848_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6139_ (.A1(\mod.pc[12] ),
    .A2(_2679_),
    .B(_2844_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6140_ (.A1(_2847_),
    .A2(_2849_),
    .B(_2850_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6141_ (.I(_2670_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_2826_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6143_ (.A1(\mod.pc_1[13] ),
    .A2(_2852_),
    .B(_2844_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6144_ (.A1(_2818_),
    .A2(_2851_),
    .B(_2853_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6145_ (.I(\mod.instr[0] ),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6146_ (.I(_2673_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6147_ (.I(_2855_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6148_ (.A1(\mod.des.des_dout[0] ),
    .A2(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6149_ (.I(_1856_),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_2858_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6151_ (.A1(_2854_),
    .A2(_2675_),
    .B1(_2857_),
    .B2(_2859_),
    .C(_2823_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6152_ (.I(\mod.instr[1] ),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6153_ (.A1(\mod.des.des_dout[1] ),
    .A2(_2856_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6154_ (.A1(_2860_),
    .A2(_2675_),
    .B1(_2861_),
    .B2(_2859_),
    .C(_2823_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6155_ (.I(\mod.instr[2] ),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6156_ (.I(_2855_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6157_ (.A1(\mod.des.des_dout[2] ),
    .A2(_2863_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6158_ (.A1(_2862_),
    .A2(_2675_),
    .B1(_2864_),
    .B2(_2859_),
    .C(_2823_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6159_ (.I(\mod.instr[3] ),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6160_ (.I(_2673_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(_2866_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6162_ (.A1(\mod.des.des_dout[3] ),
    .A2(_2863_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_2683_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6164_ (.A1(_2865_),
    .A2(_2867_),
    .B1(_2868_),
    .B2(_2859_),
    .C(_2869_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6165_ (.I(\mod.instr[4] ),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6166_ (.A1(\mod.des.des_dout[4] ),
    .A2(_2863_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6167_ (.I(_2858_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6168_ (.A1(_2870_),
    .A2(_2867_),
    .B1(_2871_),
    .B2(_2872_),
    .C(_2869_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6169_ (.I(\mod.instr[5] ),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6170_ (.A1(\mod.des.des_dout[5] ),
    .A2(_2863_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6171_ (.A1(_2873_),
    .A2(_2867_),
    .B1(_2874_),
    .B2(_2872_),
    .C(_2869_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6172_ (.I(\mod.instr[6] ),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6173_ (.I(_2855_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6174_ (.A1(\mod.des.des_dout[6] ),
    .A2(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6175_ (.A1(_2875_),
    .A2(_2867_),
    .B1(_2877_),
    .B2(_2872_),
    .C(_2869_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6176_ (.I(\mod.instr[7] ),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6177_ (.I(_2674_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6178_ (.A1(\mod.des.des_dout[7] ),
    .A2(_2876_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6179_ (.I(_2683_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6180_ (.A1(_2878_),
    .A2(_2879_),
    .B1(_2880_),
    .B2(_2872_),
    .C(_2881_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6181_ (.I(\mod.instr[8] ),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6182_ (.A1(\mod.des.des_dout[8] ),
    .A2(_2876_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6183_ (.I(_2858_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6184_ (.A1(_2882_),
    .A2(_2879_),
    .B1(_2883_),
    .B2(_2884_),
    .C(_2881_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6185_ (.I(\mod.instr[9] ),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6186_ (.A1(\mod.des.des_dout[9] ),
    .A2(_2876_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6187_ (.A1(_2885_),
    .A2(_2879_),
    .B1(_2886_),
    .B2(_2884_),
    .C(_2881_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6188_ (.I(\mod.instr[10] ),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6189_ (.I(_2855_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6190_ (.A1(\mod.des.des_dout[10] ),
    .A2(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6191_ (.A1(_2887_),
    .A2(_2879_),
    .B1(_2889_),
    .B2(_2884_),
    .C(_2881_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6192_ (.I(\mod.instr[11] ),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6193_ (.I(_2674_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6194_ (.A1(\mod.des.des_dout[11] ),
    .A2(_2888_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6195_ (.I(_2718_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6196_ (.A1(_2890_),
    .A2(_2891_),
    .B1(_2892_),
    .B2(_2884_),
    .C(_2893_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6197_ (.I(\mod.instr[12] ),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6198_ (.A1(\mod.des.des_dout[12] ),
    .A2(_2888_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6199_ (.I(_1856_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6200_ (.A1(_2894_),
    .A2(_2891_),
    .B1(_2895_),
    .B2(_2896_),
    .C(_2893_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6201_ (.I(\mod.instr[13] ),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6202_ (.A1(\mod.des.des_dout[13] ),
    .A2(_2888_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6203_ (.A1(_2897_),
    .A2(_2891_),
    .B1(_2898_),
    .B2(_2896_),
    .C(_2893_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6204_ (.I(\mod.instr[14] ),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6205_ (.I(_2673_),
    .Z(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6206_ (.A1(\mod.des.des_dout[14] ),
    .A2(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6207_ (.A1(_2899_),
    .A2(_2891_),
    .B1(_2901_),
    .B2(_2896_),
    .C(_2893_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6208_ (.I(\mod.instr[15] ),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6209_ (.I(_2674_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6210_ (.A1(\mod.des.des_dout[15] ),
    .A2(_2900_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6211_ (.I(_2718_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6212_ (.A1(_2902_),
    .A2(_2903_),
    .B1(_2904_),
    .B2(_2896_),
    .C(_2905_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6213_ (.I(\mod.instr[16] ),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6214_ (.A1(\mod.des.des_dout[16] ),
    .A2(_2900_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6215_ (.I(_1856_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6216_ (.A1(_2906_),
    .A2(_2903_),
    .B1(_2907_),
    .B2(_2908_),
    .C(_2905_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6217_ (.I(\mod.instr[17] ),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6218_ (.A1(\mod.des.des_dout[17] ),
    .A2(_2900_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6219_ (.A1(_2909_),
    .A2(_2903_),
    .B1(_2910_),
    .B2(_2908_),
    .C(_2905_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6220_ (.I(\mod.instr[18] ),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6221_ (.A1(\mod.des.des_dout[18] ),
    .A2(_2866_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6222_ (.A1(_2911_),
    .A2(_2903_),
    .B1(_2912_),
    .B2(_2908_),
    .C(_2905_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6223_ (.I(\mod.instr[19] ),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6224_ (.A1(\mod.des.des_dout[19] ),
    .A2(_2866_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6225_ (.I(_2665_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6226_ (.A1(_2913_),
    .A2(_2856_),
    .B1(_2914_),
    .B2(_2908_),
    .C(_2915_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6227_ (.I(\mod.instr[20] ),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6228_ (.A1(\mod.des.des_dout[20] ),
    .A2(_2866_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6229_ (.A1(_2916_),
    .A2(_2856_),
    .B1(_2917_),
    .B2(_2858_),
    .C(_2915_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6230_ (.A1(_2668_),
    .A2(_2681_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6231_ (.I(_2918_),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_2678_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_1346_),
    .A2(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6234_ (.A1(_2919_),
    .A2(_2921_),
    .B(_2799_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6235_ (.I(_2915_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6236_ (.A1(_3196_),
    .A2(_2671_),
    .B1(_2919_),
    .B2(\mod.instr[0] ),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6237_ (.A1(_2922_),
    .A2(_2923_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6238_ (.I(_2670_),
    .Z(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6239_ (.A1(_1750_),
    .A2(_2924_),
    .B1(_2919_),
    .B2(\mod.instr[1] ),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6240_ (.A1(_2922_),
    .A2(_2925_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6241_ (.A1(_3194_),
    .A2(_2924_),
    .B1(_2919_),
    .B2(\mod.instr[2] ),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6242_ (.A1(_2922_),
    .A2(_2926_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6243_ (.I(_2918_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6244_ (.I(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6245_ (.A1(_1817_),
    .A2(_2924_),
    .B1(_2928_),
    .B2(\mod.instr[3] ),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6246_ (.A1(_2922_),
    .A2(_2929_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6247_ (.I(_2915_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6248_ (.A1(_1816_),
    .A2(_2924_),
    .B1(_2928_),
    .B2(\mod.instr[4] ),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6249_ (.A1(_2930_),
    .A2(_2931_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6250_ (.I(_1831_),
    .Z(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6251_ (.I(_2932_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6252_ (.I(_2669_),
    .Z(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6253_ (.I(_2934_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6254_ (.A1(_2933_),
    .A2(_2935_),
    .B1(_2928_),
    .B2(\mod.instr[5] ),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6255_ (.A1(_2930_),
    .A2(_2936_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6256_ (.A1(\mod.instr_2[6] ),
    .A2(_2935_),
    .B1(_2928_),
    .B2(\mod.instr[6] ),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6257_ (.A1(_2930_),
    .A2(_2937_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6258_ (.I(_2927_),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6259_ (.A1(_1518_),
    .A2(_2935_),
    .B1(_2938_),
    .B2(\mod.instr[7] ),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6260_ (.A1(_2930_),
    .A2(_2939_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_2665_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6262_ (.I(_2940_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6263_ (.A1(_1348_),
    .A2(_2935_),
    .B1(_2938_),
    .B2(\mod.instr[8] ),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6264_ (.A1(_2941_),
    .A2(_2942_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6265_ (.I(_2934_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6266_ (.A1(_1347_),
    .A2(_2943_),
    .B1(_2938_),
    .B2(\mod.instr[9] ),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6267_ (.A1(_2941_),
    .A2(_2944_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6268_ (.A1(_1801_),
    .A2(_2943_),
    .B1(_2938_),
    .B2(\mod.instr[10] ),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6269_ (.A1(_2941_),
    .A2(_2945_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6270_ (.I(_2918_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6271_ (.A1(_1802_),
    .A2(_2943_),
    .B1(_2946_),
    .B2(\mod.instr[11] ),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6272_ (.A1(_2941_),
    .A2(_2947_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6273_ (.I(_2940_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6274_ (.A1(_0607_),
    .A2(_2943_),
    .B1(_2946_),
    .B2(\mod.instr[12] ),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6275_ (.A1(_2948_),
    .A2(_2949_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6276_ (.I(_2934_),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6277_ (.A1(_0615_),
    .A2(_2950_),
    .B1(_2946_),
    .B2(\mod.instr[13] ),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6278_ (.A1(_2948_),
    .A2(_2951_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6279_ (.A1(_0445_),
    .A2(_2950_),
    .B1(_2946_),
    .B2(\mod.instr[14] ),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6280_ (.A1(_2948_),
    .A2(_2952_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6281_ (.I(_2918_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6282_ (.A1(_0585_),
    .A2(_2950_),
    .B1(_2953_),
    .B2(\mod.instr[15] ),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6283_ (.A1(_2948_),
    .A2(_2954_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6284_ (.I(_2940_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6285_ (.A1(_0697_),
    .A2(_2950_),
    .B1(_2953_),
    .B2(\mod.instr[16] ),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6286_ (.A1(_2955_),
    .A2(_2956_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6287_ (.I(_2934_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6288_ (.A1(_0476_),
    .A2(_2957_),
    .B1(_2953_),
    .B2(\mod.instr[17] ),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6289_ (.A1(_2955_),
    .A2(_2958_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6290_ (.A1(\mod.funct7[0] ),
    .A2(_2957_),
    .B1(_2953_),
    .B2(\mod.instr[18] ),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6291_ (.A1(_2955_),
    .A2(_2959_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6292_ (.A1(\mod.funct7[1] ),
    .A2(_2957_),
    .B1(_2927_),
    .B2(\mod.instr[19] ),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6293_ (.A1(_2955_),
    .A2(_2960_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6294_ (.I(_2940_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6295_ (.A1(_1177_),
    .A2(_2957_),
    .B1(_2927_),
    .B2(\mod.instr[20] ),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6296_ (.A1(_2961_),
    .A2(_2962_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6297_ (.I(_2096_),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6298_ (.I(_2963_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6299_ (.A1(\mod.pc_1[0] ),
    .A2(_2679_),
    .B(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6300_ (.A1(_3224_),
    .A2(_2849_),
    .B(_2965_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_2678_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6302_ (.A1(\mod.pc_1[1] ),
    .A2(_2966_),
    .B(_2964_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6303_ (.A1(_0830_),
    .A2(_2849_),
    .B(_2967_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6304_ (.A1(\mod.pc_1[2] ),
    .A2(_2966_),
    .B(_2964_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6305_ (.A1(_0813_),
    .A2(_2849_),
    .B(_2968_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6306_ (.I(_2848_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6307_ (.A1(\mod.pc_1[3] ),
    .A2(_2966_),
    .B(_2964_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6308_ (.A1(_0799_),
    .A2(_2969_),
    .B(_2970_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6309_ (.I(_2963_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6310_ (.A1(\mod.pc_1[4] ),
    .A2(_2966_),
    .B(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6311_ (.A1(_2161_),
    .A2(_2969_),
    .B(_2972_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6312_ (.I(_2677_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6313_ (.A1(\mod.pc_1[5] ),
    .A2(_2973_),
    .B(_2971_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6314_ (.A1(_0769_),
    .A2(_2969_),
    .B(_2974_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6315_ (.I(_1968_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6316_ (.A1(\mod.pc_1[6] ),
    .A2(_2973_),
    .B(_2971_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6317_ (.A1(_2975_),
    .A2(_2969_),
    .B(_2976_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6318_ (.I(_2678_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6319_ (.A1(\mod.pc_1[7] ),
    .A2(_2973_),
    .B(_2971_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6320_ (.A1(_0740_),
    .A2(_2977_),
    .B(_2978_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6321_ (.I(_2963_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6322_ (.A1(\mod.pc_1[8] ),
    .A2(_2973_),
    .B(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6323_ (.A1(_1092_),
    .A2(_2977_),
    .B(_2980_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6324_ (.I(_2024_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6325_ (.I(_2677_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6326_ (.A1(\mod.pc_1[9] ),
    .A2(_2982_),
    .B(_2979_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6327_ (.A1(_2981_),
    .A2(_2977_),
    .B(_2983_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6328_ (.A1(\mod.pc_1[10] ),
    .A2(_2982_),
    .B(_2979_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6329_ (.A1(_2043_),
    .A2(_2977_),
    .B(_2984_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6330_ (.I(_2057_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6331_ (.A1(\mod.pc_1[11] ),
    .A2(_2982_),
    .B(_2979_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6332_ (.A1(_2985_),
    .A2(_2920_),
    .B(_2986_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6333_ (.I(_2963_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6334_ (.A1(\mod.pc_1[12] ),
    .A2(_2982_),
    .B(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6335_ (.A1(_1138_),
    .A2(_2920_),
    .B(_2988_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6336_ (.A1(\mod.pc_1[13] ),
    .A2(_2848_),
    .B(_2987_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6337_ (.A1(_1209_),
    .A2(_2920_),
    .B(_2989_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6338_ (.A1(\mod.valid_out3 ),
    .A2(_2112_),
    .A3(_2848_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6339_ (.A1(_2111_),
    .A2(_2990_),
    .B(_2799_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6340_ (.A1(_0851_),
    .A2(_1760_),
    .A3(_2668_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6341_ (.I(_2991_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6342_ (.A1(_3214_),
    .A2(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6343_ (.A1(net20),
    .A2(_2111_),
    .B1(_2993_),
    .B2(_1346_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6344_ (.A1(_2961_),
    .A2(_2994_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6345_ (.A1(\mod.ri_3 ),
    .A2(_2852_),
    .B(_2987_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6346_ (.A1(_0914_),
    .A2(_2851_),
    .B(_2995_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6347_ (.A1(\mod.ins_ldr_3 ),
    .A2(_2679_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6348_ (.A1(_2992_),
    .A2(_2996_),
    .B(_2799_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6349_ (.A1(\mod.rd_3[0] ),
    .A2(_2852_),
    .B(_2987_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6350_ (.A1(_1818_),
    .A2(_2851_),
    .B(_2997_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6351_ (.A1(\mod.rd_3[1] ),
    .A2(_2852_),
    .B(_2097_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6352_ (.A1(_1821_),
    .A2(_2851_),
    .B(_2998_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6353_ (.I(_2098_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6354_ (.A1(\mod.rd_3[2] ),
    .A2(_2824_),
    .B(_2097_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6355_ (.A1(_2999_),
    .A2(_2671_),
    .B(_3000_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6356_ (.A1(\mod.rd_3[3] ),
    .A2(_2824_),
    .B(_2097_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6357_ (.A1(_2104_),
    .A2(_2671_),
    .B(_3001_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6358_ (.A1(_2698_),
    .A2(_1763_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6359_ (.I(_3002_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6360_ (.A1(_1782_),
    .A2(_0003_),
    .A3(_3003_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6361_ (.I(_3004_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6362_ (.A1(_1781_),
    .A2(_3003_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6363_ (.I(_1820_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6364_ (.A1(\mod.instr_2[6] ),
    .A2(_2991_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6365_ (.I(_3007_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6366_ (.A1(_2999_),
    .A2(_3006_),
    .A3(_3008_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6367_ (.I(_2666_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6368_ (.A1(_3005_),
    .A2(_3009_),
    .B(_3010_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6369_ (.A1(_1780_),
    .A2(_3003_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6370_ (.I(_1826_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6371_ (.A1(_2999_),
    .A2(_3012_),
    .A3(_3008_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6372_ (.A1(_3011_),
    .A2(_3013_),
    .B(_3010_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_1779_),
    .A2(_3003_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6374_ (.I(_1823_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6375_ (.A1(_2999_),
    .A2(_3015_),
    .A3(_3008_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6376_ (.A1(_3014_),
    .A2(_3016_),
    .B(_3010_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6377_ (.I(_3002_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6378_ (.A1(_1767_),
    .A2(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6379_ (.A1(_2933_),
    .A2(_1828_),
    .A3(_3008_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6380_ (.A1(_3018_),
    .A2(_3019_),
    .B(_3010_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6381_ (.A1(_1766_),
    .A2(_3017_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6382_ (.A1(_2933_),
    .A2(_3006_),
    .A3(_3007_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6383_ (.I(_2666_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6384_ (.A1(_3020_),
    .A2(_3021_),
    .B(_3022_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6385_ (.A1(_1765_),
    .A2(_3017_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6386_ (.A1(_2933_),
    .A2(_3012_),
    .A3(_3007_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6387_ (.A1(_3023_),
    .A2(_3024_),
    .B(_3022_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6388_ (.A1(_1764_),
    .A2(_3017_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6389_ (.I(_2932_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6390_ (.A1(_3026_),
    .A2(_3015_),
    .A3(_3007_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6391_ (.A1(_3025_),
    .A2(_3027_),
    .B(_3022_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6392_ (.I(_3002_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6393_ (.A1(_2104_),
    .A2(_2932_),
    .A3(_2992_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6394_ (.A1(_1772_),
    .A2(_3028_),
    .B1(_3029_),
    .B2(_1828_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6395_ (.A1(_2961_),
    .A2(_3030_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6396_ (.A1(_1771_),
    .A2(_3028_),
    .B1(_3029_),
    .B2(_3006_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_2961_),
    .A2(_3031_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6398_ (.A1(_1770_),
    .A2(_3028_),
    .B1(_3029_),
    .B2(_3012_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6399_ (.A1(_2684_),
    .A2(_3032_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6400_ (.A1(_1769_),
    .A2(_3028_),
    .B1(_3029_),
    .B2(_3015_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6401_ (.A1(_2684_),
    .A2(_3033_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6402_ (.I(_3002_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6403_ (.A1(_1777_),
    .A2(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6404_ (.A1(_2104_),
    .A2(_2992_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6405_ (.A1(_3026_),
    .A2(_1828_),
    .A3(_3036_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6406_ (.A1(_3035_),
    .A2(_3037_),
    .B(_3022_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(_1776_),
    .A2(_3034_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6408_ (.A1(_3026_),
    .A2(_3006_),
    .A3(_3036_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6409_ (.A1(_3038_),
    .A2(_3039_),
    .B(_2732_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6410_ (.A1(_1775_),
    .A2(_3034_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6411_ (.A1(_3026_),
    .A2(_3012_),
    .A3(_3036_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6412_ (.A1(_3040_),
    .A2(_3041_),
    .B(_2732_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6413_ (.A1(_1774_),
    .A2(_3034_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6414_ (.A1(_2932_),
    .A2(_3015_),
    .A3(_3036_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6415_ (.A1(_3042_),
    .A2(_3043_),
    .B(_2732_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6416_ (.A1(\mod.des.des_counter[0] ),
    .A2(\mod.des.des_counter[1] ),
    .A3(\mod.des.des_counter[2] ),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6417_ (.I(_3044_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6418_ (.I0(\mod.des.des_dout[0] ),
    .I1(net16),
    .S(_3045_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6419_ (.I(_3046_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6420_ (.I0(\mod.des.des_dout[1] ),
    .I1(net17),
    .S(_3045_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6421_ (.I(_3047_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6422_ (.I0(\mod.des.des_dout[2] ),
    .I1(net18),
    .S(_3045_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6423_ (.I(_3048_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6424_ (.I0(\mod.des.des_dout[3] ),
    .I1(net19),
    .S(_3045_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6425_ (.I(_3049_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6426_ (.I(_3044_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6427_ (.I0(\mod.des.des_dout[4] ),
    .I1(net2),
    .S(_3050_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6428_ (.I(_3051_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6429_ (.I0(\mod.des.des_dout[5] ),
    .I1(net3),
    .S(_3050_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6430_ (.I(_3052_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6431_ (.I0(\mod.des.des_dout[6] ),
    .I1(net4),
    .S(_3050_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6432_ (.I(_3053_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6433_ (.I0(\mod.des.des_dout[7] ),
    .I1(net5),
    .S(_3050_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6434_ (.I(_3054_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6435_ (.I(_3044_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6436_ (.I0(\mod.des.des_dout[8] ),
    .I1(net6),
    .S(_3055_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6437_ (.I(_3056_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6438_ (.I0(\mod.des.des_dout[9] ),
    .I1(net7),
    .S(_3055_),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_3057_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6440_ (.I0(\mod.des.des_dout[10] ),
    .I1(net8),
    .S(_3055_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_3058_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6442_ (.I0(\mod.des.des_dout[11] ),
    .I1(net9),
    .S(_3055_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_3059_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6444_ (.I0(\mod.des.des_dout[12] ),
    .I1(net10),
    .S(_3044_),
    .Z(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6445_ (.I(_3060_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_2286_),
    .A2(_2583_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6447_ (.I(_3061_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6448_ (.I(_3062_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6449_ (.I(_3061_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6450_ (.I(_3064_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6451_ (.A1(\mod.registers.r15[0] ),
    .A2(_3065_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6452_ (.A1(_2344_),
    .A2(_3063_),
    .B(_3066_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6453_ (.A1(\mod.registers.r15[1] ),
    .A2(_3065_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6454_ (.A1(_2352_),
    .A2(_3063_),
    .B(_3067_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6455_ (.A1(\mod.registers.r15[2] ),
    .A2(_3065_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6456_ (.A1(_2355_),
    .A2(_3063_),
    .B(_3068_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6457_ (.A1(\mod.registers.r15[3] ),
    .A2(_3065_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6458_ (.A1(_2358_),
    .A2(_3063_),
    .B(_3069_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6459_ (.I(_3062_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6460_ (.I(_3064_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6461_ (.A1(\mod.registers.r15[4] ),
    .A2(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6462_ (.A1(_2361_),
    .A2(_3070_),
    .B(_3072_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6463_ (.A1(\mod.registers.r15[5] ),
    .A2(_3071_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6464_ (.A1(_2366_),
    .A2(_3070_),
    .B(_3073_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6465_ (.A1(\mod.registers.r15[6] ),
    .A2(_3071_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6466_ (.A1(_2369_),
    .A2(_3070_),
    .B(_3074_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6467_ (.A1(\mod.registers.r15[7] ),
    .A2(_3071_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6468_ (.A1(_2372_),
    .A2(_3070_),
    .B(_3075_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6469_ (.I(_3062_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6470_ (.I(_3064_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6471_ (.A1(\mod.registers.r15[8] ),
    .A2(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6472_ (.A1(_2375_),
    .A2(_3076_),
    .B(_3078_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(\mod.registers.r15[9] ),
    .A2(_3077_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6474_ (.A1(_2380_),
    .A2(_3076_),
    .B(_3079_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(\mod.registers.r15[10] ),
    .A2(_3077_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6476_ (.A1(_2383_),
    .A2(_3076_),
    .B(_3080_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6477_ (.A1(\mod.registers.r15[11] ),
    .A2(_3077_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6478_ (.A1(_2386_),
    .A2(_3076_),
    .B(_3081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6479_ (.I(_3062_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6480_ (.I(_3064_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6481_ (.A1(\mod.registers.r15[12] ),
    .A2(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6482_ (.A1(_2389_),
    .A2(_3082_),
    .B(_3084_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6483_ (.A1(\mod.registers.r15[13] ),
    .A2(_3083_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6484_ (.A1(_2394_),
    .A2(_3082_),
    .B(_3085_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6485_ (.A1(\mod.registers.r15[14] ),
    .A2(_3083_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6486_ (.A1(_2397_),
    .A2(_3082_),
    .B(_3086_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6487_ (.A1(\mod.registers.r15[15] ),
    .A2(_3083_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6488_ (.A1(_2400_),
    .A2(_3082_),
    .B(_3087_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6489_ (.A1(\mod.des.des_counter[2] ),
    .A2(_1872_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6490_ (.I(_3088_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6491_ (.I0(\mod.des.des_dout[13] ),
    .I1(net16),
    .S(_3089_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6492_ (.I(_3090_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6493_ (.I0(\mod.des.des_dout[14] ),
    .I1(net17),
    .S(_3089_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6494_ (.I(_3091_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6495_ (.I0(\mod.des.des_dout[15] ),
    .I1(net18),
    .S(_3089_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6496_ (.I(_3092_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6497_ (.I0(\mod.des.des_dout[16] ),
    .I1(net19),
    .S(_3089_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6498_ (.I(_3093_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6499_ (.I(_3088_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6500_ (.I0(\mod.des.des_dout[17] ),
    .I1(net2),
    .S(_3094_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6501_ (.I(_3095_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6502_ (.I0(\mod.des.des_dout[18] ),
    .I1(net3),
    .S(_3094_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6503_ (.I(_3096_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6504_ (.I0(\mod.des.des_dout[19] ),
    .I1(net4),
    .S(_3094_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6505_ (.I(_3097_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6506_ (.I0(\mod.des.des_dout[20] ),
    .I1(net5),
    .S(_3094_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6507_ (.I(_3098_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6508_ (.I(_3088_),
    .Z(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6509_ (.I0(\mod.des.des_dout[21] ),
    .I1(net6),
    .S(_3099_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6510_ (.I(_3100_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6511_ (.I0(\mod.des.des_dout[22] ),
    .I1(net7),
    .S(_3099_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6512_ (.I(_3101_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6513_ (.I0(\mod.des.des_dout[23] ),
    .I1(net8),
    .S(_3099_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6514_ (.I(_3102_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6515_ (.I0(\mod.des.des_dout[24] ),
    .I1(net9),
    .S(_3099_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6516_ (.I(_3103_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6517_ (.I0(\mod.des.des_dout[25] ),
    .I1(net10),
    .S(_3088_),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6518_ (.I(_3104_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6519_ (.A1(\mod.des.des_counter[2] ),
    .A2(_1945_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6520_ (.I(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6521_ (.I(_3106_),
    .Z(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6522_ (.I0(net16),
    .I1(\mod.des.des_dout[26] ),
    .S(_3107_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6523_ (.I(_3108_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6524_ (.I0(net17),
    .I1(\mod.des.des_dout[27] ),
    .S(_3107_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6525_ (.I(_3109_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6526_ (.I0(net18),
    .I1(\mod.des.des_dout[28] ),
    .S(_3107_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6527_ (.I(_3110_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6528_ (.I0(net19),
    .I1(\mod.des.des_dout[29] ),
    .S(_3107_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_3111_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6530_ (.I(_3105_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6531_ (.I0(net2),
    .I1(\mod.des.des_dout[30] ),
    .S(_3112_),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6532_ (.I(_3113_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6533_ (.I0(net3),
    .I1(\mod.des.des_dout[31] ),
    .S(_3112_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6534_ (.I(_3114_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6535_ (.I0(net4),
    .I1(\mod.des.des_dout[32] ),
    .S(_3112_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6536_ (.I(_3115_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6537_ (.I0(net5),
    .I1(\mod.des.des_dout[33] ),
    .S(_3112_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6538_ (.I(_3116_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6539_ (.I0(net6),
    .I1(\mod.des.des_dout[34] ),
    .S(_3106_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6540_ (.I(_3117_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6541_ (.I0(net7),
    .I1(\mod.des.des_dout[35] ),
    .S(_3106_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6542_ (.I(_3118_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6543_ (.I0(net8),
    .I1(\mod.des.des_dout[36] ),
    .S(_3106_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6544_ (.I(_3119_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6545_ (.D(_0111_),
    .RN(_0003_),
    .CLK(net206),
    .Q(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6546_ (.D(_0112_),
    .CLK(net140),
    .Q(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6547_ (.D(_0113_),
    .CLK(net137),
    .Q(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6548_ (.D(_0114_),
    .CLK(net137),
    .Q(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6549_ (.D(_0115_),
    .CLK(net139),
    .Q(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6550_ (.D(_0116_),
    .CLK(net130),
    .Q(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6551_ (.D(_0117_),
    .CLK(net129),
    .Q(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6552_ (.D(_0118_),
    .CLK(net141),
    .Q(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6553_ (.D(_0119_),
    .CLK(net133),
    .Q(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6554_ (.D(_0120_),
    .CLK(net82),
    .Q(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6555_ (.D(_0121_),
    .CLK(net85),
    .Q(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6556_ (.D(_0122_),
    .CLK(net82),
    .Q(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6557_ (.D(_0123_),
    .CLK(net85),
    .Q(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6558_ (.D(_0124_),
    .CLK(net78),
    .Q(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6559_ (.D(_0125_),
    .CLK(net74),
    .Q(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6560_ (.D(_0126_),
    .CLK(net74),
    .Q(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6561_ (.D(_0127_),
    .CLK(net78),
    .Q(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6562_ (.D(_0128_),
    .CLK(net134),
    .Q(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6563_ (.D(_0129_),
    .CLK(net138),
    .Q(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6564_ (.D(_0130_),
    .CLK(net134),
    .Q(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6565_ (.D(_0131_),
    .CLK(net138),
    .Q(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6566_ (.D(_0132_),
    .CLK(net130),
    .Q(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6567_ (.D(_0133_),
    .CLK(net129),
    .Q(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6568_ (.D(_0134_),
    .CLK(net129),
    .Q(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6569_ (.D(_0135_),
    .CLK(net129),
    .Q(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6570_ (.D(_0136_),
    .CLK(net80),
    .Q(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6571_ (.D(_0137_),
    .CLK(net86),
    .Q(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6572_ (.D(_0138_),
    .CLK(net128),
    .Q(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6573_ (.D(_0139_),
    .CLK(net82),
    .Q(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6574_ (.D(_0140_),
    .CLK(net76),
    .Q(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6575_ (.D(_0141_),
    .CLK(net75),
    .Q(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6576_ (.D(_0142_),
    .CLK(net76),
    .Q(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6577_ (.D(_0143_),
    .CLK(net75),
    .Q(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6578_ (.D(_0144_),
    .CLK(net133),
    .Q(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6579_ (.D(_0145_),
    .CLK(net137),
    .Q(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6580_ (.D(_0146_),
    .CLK(net133),
    .Q(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6581_ (.D(_0147_),
    .CLK(net137),
    .Q(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6582_ (.D(_0148_),
    .CLK(net128),
    .Q(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6583_ (.D(_0149_),
    .CLK(net128),
    .Q(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6584_ (.D(_0150_),
    .CLK(net127),
    .Q(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6585_ (.D(_0151_),
    .CLK(net128),
    .Q(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6586_ (.D(_0152_),
    .CLK(net80),
    .Q(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6587_ (.D(_0153_),
    .CLK(net81),
    .Q(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6588_ (.D(_0154_),
    .CLK(net81),
    .Q(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6589_ (.D(_0155_),
    .CLK(net81),
    .Q(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6590_ (.D(_0156_),
    .CLK(net43),
    .Q(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6591_ (.D(_0157_),
    .CLK(net74),
    .Q(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6592_ (.D(_0158_),
    .CLK(net74),
    .Q(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6593_ (.D(_0159_),
    .CLK(net75),
    .Q(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6594_ (.D(_0160_),
    .CLK(net140),
    .Q(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6595_ (.D(_0161_),
    .CLK(net138),
    .Q(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6596_ (.D(_0162_),
    .CLK(net138),
    .Q(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6597_ (.D(_0163_),
    .CLK(net139),
    .Q(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6598_ (.D(_0164_),
    .CLK(net126),
    .Q(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6599_ (.D(_0165_),
    .CLK(net126),
    .Q(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6600_ (.D(_0166_),
    .CLK(net127),
    .Q(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6601_ (.D(_0167_),
    .CLK(net126),
    .Q(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6602_ (.D(_0168_),
    .CLK(net83),
    .Q(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6603_ (.D(_0169_),
    .CLK(net82),
    .Q(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6604_ (.D(_0170_),
    .CLK(net126),
    .Q(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6605_ (.D(_0171_),
    .CLK(net83),
    .Q(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6606_ (.D(_0172_),
    .CLK(net77),
    .Q(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6607_ (.D(_0173_),
    .CLK(net77),
    .Q(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6608_ (.D(_0174_),
    .CLK(net79),
    .Q(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6609_ (.D(_0175_),
    .CLK(net79),
    .Q(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6610_ (.D(_0176_),
    .CLK(net110),
    .Q(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6611_ (.D(_0177_),
    .CLK(net110),
    .Q(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6612_ (.D(_0178_),
    .CLK(net94),
    .Q(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6613_ (.D(_0179_),
    .CLK(net110),
    .Q(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6614_ (.D(_0180_),
    .CLK(net95),
    .Q(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6615_ (.D(_0181_),
    .CLK(net94),
    .Q(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6616_ (.D(_0182_),
    .CLK(net94),
    .Q(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6617_ (.D(_0183_),
    .CLK(net89),
    .Q(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6618_ (.D(_0184_),
    .CLK(net56),
    .Q(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6619_ (.D(_0185_),
    .CLK(net52),
    .Q(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6620_ (.D(_0186_),
    .CLK(net90),
    .Q(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6621_ (.D(_0187_),
    .CLK(net58),
    .Q(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6622_ (.D(_0188_),
    .CLK(net51),
    .Q(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6623_ (.D(_0189_),
    .CLK(net51),
    .Q(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6624_ (.D(_0190_),
    .CLK(net38),
    .Q(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6625_ (.D(_0191_),
    .CLK(net40),
    .Q(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6626_ (.D(_0192_),
    .CLK(net112),
    .Q(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6627_ (.D(_0193_),
    .CLK(net110),
    .Q(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6628_ (.D(_0194_),
    .CLK(net98),
    .Q(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6629_ (.D(_0195_),
    .CLK(net113),
    .Q(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6630_ (.D(_0196_),
    .CLK(net89),
    .Q(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6631_ (.D(_0197_),
    .CLK(net90),
    .Q(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6632_ (.D(_0198_),
    .CLK(net95),
    .Q(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6633_ (.D(_0199_),
    .CLK(net89),
    .Q(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6634_ (.D(_0200_),
    .CLK(net57),
    .Q(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6635_ (.D(_0201_),
    .CLK(net56),
    .Q(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6636_ (.D(_0202_),
    .CLK(net57),
    .Q(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6637_ (.D(_0203_),
    .CLK(net56),
    .Q(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6638_ (.D(_0204_),
    .CLK(net51),
    .Q(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6639_ (.D(_0205_),
    .CLK(net51),
    .Q(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6640_ (.D(_0206_),
    .CLK(net40),
    .Q(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6641_ (.D(_0207_),
    .CLK(net40),
    .Q(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6642_ (.D(_0208_),
    .CLK(net111),
    .Q(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6643_ (.D(_0209_),
    .CLK(net111),
    .Q(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6644_ (.D(_0210_),
    .CLK(net97),
    .Q(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6645_ (.D(_0211_),
    .CLK(net111),
    .Q(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6646_ (.D(_0212_),
    .CLK(net89),
    .Q(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6647_ (.D(_0213_),
    .CLK(net95),
    .Q(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6648_ (.D(_0214_),
    .CLK(net94),
    .Q(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6649_ (.D(_0215_),
    .CLK(net93),
    .Q(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6650_ (.D(_0216_),
    .CLK(net57),
    .Q(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6651_ (.D(_0217_),
    .CLK(net56),
    .Q(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6652_ (.D(_0218_),
    .CLK(net90),
    .Q(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6653_ (.D(_0219_),
    .CLK(net52),
    .Q(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6654_ (.D(_0220_),
    .CLK(net53),
    .Q(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6655_ (.D(_0221_),
    .CLK(net53),
    .Q(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6656_ (.D(_0222_),
    .CLK(net39),
    .Q(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6657_ (.D(_0223_),
    .CLK(net38),
    .Q(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6658_ (.D(_0224_),
    .CLK(net112),
    .Q(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6659_ (.D(_0225_),
    .CLK(net115),
    .Q(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6660_ (.D(_0226_),
    .CLK(net97),
    .Q(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6661_ (.D(_0227_),
    .CLK(net111),
    .Q(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6662_ (.D(_0228_),
    .CLK(net96),
    .Q(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6663_ (.D(_0229_),
    .CLK(net91),
    .Q(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6664_ (.D(_0230_),
    .CLK(net96),
    .Q(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6665_ (.D(_0231_),
    .CLK(net92),
    .Q(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6666_ (.D(_0232_),
    .CLK(net59),
    .Q(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6667_ (.D(_0233_),
    .CLK(net58),
    .Q(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6668_ (.D(_0234_),
    .CLK(net91),
    .Q(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6669_ (.D(_0235_),
    .CLK(net58),
    .Q(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6670_ (.D(_0236_),
    .CLK(net53),
    .Q(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6671_ (.D(_0237_),
    .CLK(net53),
    .Q(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6672_ (.D(_0238_),
    .CLK(net38),
    .Q(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6673_ (.D(_0239_),
    .CLK(net38),
    .Q(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6674_ (.D(_0240_),
    .CLK(net132),
    .Q(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6675_ (.D(_0241_),
    .CLK(net132),
    .Q(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6676_ (.D(_0242_),
    .CLK(net121),
    .Q(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6677_ (.D(_0243_),
    .CLK(net131),
    .Q(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6678_ (.D(_0244_),
    .CLK(net105),
    .Q(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6679_ (.D(_0245_),
    .CLK(net101),
    .Q(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6680_ (.D(_0246_),
    .CLK(net105),
    .Q(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6681_ (.D(_0247_),
    .CLK(net102),
    .Q(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6682_ (.D(_0248_),
    .CLK(net80),
    .Q(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6683_ (.D(_0249_),
    .CLK(net68),
    .Q(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6684_ (.D(_0250_),
    .CLK(net69),
    .Q(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6685_ (.D(_0251_),
    .CLK(net64),
    .Q(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6686_ (.D(_0252_),
    .CLK(net43),
    .Q(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6687_ (.D(_0253_),
    .CLK(net43),
    .Q(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6688_ (.D(_0254_),
    .CLK(net44),
    .Q(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6689_ (.D(_0255_),
    .CLK(net43),
    .Q(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6690_ (.D(_0256_),
    .CLK(net131),
    .Q(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6691_ (.D(_0257_),
    .CLK(net120),
    .Q(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6692_ (.D(_0258_),
    .CLK(net120),
    .Q(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6693_ (.D(_0259_),
    .CLK(net131),
    .Q(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6694_ (.D(_0260_),
    .CLK(net105),
    .Q(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6695_ (.D(_0261_),
    .CLK(net101),
    .Q(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6696_ (.D(_0262_),
    .CLK(net106),
    .Q(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6697_ (.D(_0263_),
    .CLK(net101),
    .Q(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6698_ (.D(_0264_),
    .CLK(net66),
    .Q(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6699_ (.D(_0265_),
    .CLK(net66),
    .Q(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6700_ (.D(_0266_),
    .CLK(net69),
    .Q(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6701_ (.D(_0267_),
    .CLK(net68),
    .Q(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6702_ (.D(_0268_),
    .CLK(net42),
    .Q(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6703_ (.D(_0269_),
    .CLK(net42),
    .Q(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6704_ (.D(_0270_),
    .CLK(net45),
    .Q(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6705_ (.D(_0271_),
    .CLK(net42),
    .Q(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6706_ (.D(_0272_),
    .CLK(net131),
    .Q(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6707_ (.D(_0273_),
    .CLK(net120),
    .Q(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6708_ (.D(_0274_),
    .CLK(net120),
    .Q(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6709_ (.D(_0275_),
    .CLK(net133),
    .Q(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6710_ (.D(_0276_),
    .CLK(net106),
    .Q(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6711_ (.D(_0277_),
    .CLK(net105),
    .Q(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6712_ (.D(_0278_),
    .CLK(net117),
    .Q(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6713_ (.D(_0279_),
    .CLK(net117),
    .Q(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6714_ (.D(_0280_),
    .CLK(net80),
    .Q(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6715_ (.D(_0281_),
    .CLK(net68),
    .Q(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6716_ (.D(_0282_),
    .CLK(net68),
    .Q(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6717_ (.D(_0283_),
    .CLK(net64),
    .Q(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6718_ (.D(_0284_),
    .CLK(net47),
    .Q(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6719_ (.D(_0285_),
    .CLK(net48),
    .Q(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6720_ (.D(_0286_),
    .CLK(net44),
    .Q(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6721_ (.D(_0287_),
    .CLK(net44),
    .Q(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6722_ (.D(_0288_),
    .CLK(net132),
    .Q(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6723_ (.D(_0289_),
    .CLK(net121),
    .Q(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6724_ (.D(_0290_),
    .CLK(net121),
    .Q(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6725_ (.D(_0291_),
    .CLK(net134),
    .Q(\mod.registers.r12[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6726_ (.D(_0292_),
    .CLK(net106),
    .Q(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6727_ (.D(_0293_),
    .CLK(net104),
    .Q(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6728_ (.D(_0294_),
    .CLK(net117),
    .Q(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6729_ (.D(_0295_),
    .CLK(net115),
    .Q(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6730_ (.D(_0296_),
    .CLK(net66),
    .Q(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6731_ (.D(_0297_),
    .CLK(net63),
    .Q(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6732_ (.D(_0298_),
    .CLK(net101),
    .Q(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6733_ (.D(_0299_),
    .CLK(net65),
    .Q(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6734_ (.D(_0300_),
    .CLK(net46),
    .Q(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6735_ (.D(_0301_),
    .CLK(net46),
    .Q(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6736_ (.D(_0302_),
    .CLK(net42),
    .Q(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6737_ (.D(_0303_),
    .CLK(net46),
    .Q(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6738_ (.D(_0304_),
    .CLK(net122),
    .Q(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6739_ (.D(_0305_),
    .CLK(net116),
    .Q(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6740_ (.D(_0306_),
    .CLK(net115),
    .Q(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6741_ (.D(_0307_),
    .CLK(net116),
    .Q(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6742_ (.D(_0308_),
    .CLK(net103),
    .Q(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6743_ (.D(_0309_),
    .CLK(net103),
    .Q(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6744_ (.D(_0310_),
    .CLK(net104),
    .Q(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6745_ (.D(_0311_),
    .CLK(net102),
    .Q(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6746_ (.D(_0312_),
    .CLK(net67),
    .Q(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6747_ (.D(_0313_),
    .CLK(net63),
    .Q(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6748_ (.D(_0314_),
    .CLK(net100),
    .Q(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6749_ (.D(_0315_),
    .CLK(net63),
    .Q(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6750_ (.D(_0316_),
    .CLK(net62),
    .Q(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6751_ (.D(_0317_),
    .CLK(net62),
    .Q(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6752_ (.D(_0318_),
    .CLK(net46),
    .Q(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6753_ (.D(_0319_),
    .CLK(net47),
    .Q(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6754_ (.D(_0320_),
    .CLK(net118),
    .Q(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6755_ (.D(_0321_),
    .CLK(net115),
    .Q(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6756_ (.D(_0322_),
    .CLK(net117),
    .Q(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6757_ (.D(_0323_),
    .CLK(net118),
    .Q(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6758_ (.D(_0324_),
    .CLK(net103),
    .Q(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6759_ (.D(_0325_),
    .CLK(net100),
    .Q(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6760_ (.D(_0326_),
    .CLK(net103),
    .Q(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6761_ (.D(_0327_),
    .CLK(net100),
    .Q(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6762_ (.D(_0328_),
    .CLK(net67),
    .Q(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6763_ (.D(_0329_),
    .CLK(net58),
    .Q(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6764_ (.D(_0330_),
    .CLK(net100),
    .Q(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6765_ (.D(_0331_),
    .CLK(net66),
    .Q(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6766_ (.D(_0332_),
    .CLK(net64),
    .Q(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6767_ (.D(_0333_),
    .CLK(net64),
    .Q(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6768_ (.D(_0334_),
    .CLK(net47),
    .Q(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6769_ (.D(_0335_),
    .CLK(net48),
    .Q(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6770_ (.D(_0000_),
    .SETN(_0004_),
    .CLK(net206),
    .Q(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6771_ (.D(_0001_),
    .SETN(_0005_),
    .CLK(net206),
    .Q(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6772_ (.D(_0002_),
    .SETN(_0006_),
    .CLK(net218),
    .Q(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6773_ (.D(_0336_),
    .CLK(net185),
    .Q(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6774_ (.D(_0337_),
    .CLK(net190),
    .Q(\mod.valid1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6775_ (.D(_0338_),
    .CLK(net163),
    .Q(\mod.pc0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6776_ (.D(_0339_),
    .CLK(net147),
    .Q(\mod.pc0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6777_ (.D(_0340_),
    .CLK(net146),
    .Q(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6778_ (.D(_0341_),
    .CLK(net146),
    .Q(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6779_ (.D(_0342_),
    .CLK(net146),
    .Q(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6780_ (.D(_0343_),
    .CLK(net150),
    .Q(\mod.pc0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6781_ (.D(_0344_),
    .CLK(net150),
    .Q(\mod.pc0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6782_ (.D(_0345_),
    .CLK(net150),
    .Q(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6783_ (.D(_0346_),
    .CLK(net147),
    .Q(\mod.pc0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6784_ (.D(_0347_),
    .CLK(net148),
    .Q(\mod.pc0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6785_ (.D(_0348_),
    .CLK(net150),
    .Q(\mod.pc0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6786_ (.D(_0349_),
    .CLK(net147),
    .Q(\mod.pc0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6787_ (.D(_0350_),
    .CLK(net149),
    .Q(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6788_ (.D(_0351_),
    .CLK(net146),
    .Q(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6789_ (.D(_0352_),
    .CLK(net157),
    .Q(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6790_ (.D(_0353_),
    .CLK(net157),
    .Q(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6791_ (.D(_0354_),
    .CLK(net155),
    .Q(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6792_ (.D(_0355_),
    .CLK(net157),
    .Q(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6793_ (.D(_0356_),
    .CLK(net149),
    .Q(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6794_ (.D(_0357_),
    .CLK(net156),
    .Q(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6795_ (.D(_0358_),
    .CLK(net155),
    .Q(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6796_ (.D(_0359_),
    .CLK(net187),
    .Q(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6797_ (.D(_0360_),
    .CLK(net149),
    .Q(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6798_ (.D(_0361_),
    .CLK(net156),
    .Q(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6799_ (.D(_0362_),
    .CLK(net155),
    .Q(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6800_ (.D(_0363_),
    .CLK(net155),
    .Q(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6801_ (.D(_0364_),
    .CLK(net162),
    .Q(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6802_ (.D(_0365_),
    .CLK(net154),
    .Q(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6803_ (.D(_0366_),
    .CLK(net158),
    .Q(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6804_ (.D(_0367_),
    .CLK(net158),
    .Q(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6805_ (.D(_0368_),
    .CLK(net190),
    .Q(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6806_ (.D(_0369_),
    .CLK(net157),
    .Q(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6807_ (.D(_0370_),
    .CLK(net189),
    .Q(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6808_ (.D(_0371_),
    .CLK(net189),
    .Q(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6809_ (.D(_0372_),
    .CLK(net188),
    .Q(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6810_ (.D(_0373_),
    .CLK(net187),
    .Q(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6811_ (.D(_0374_),
    .CLK(net159),
    .Q(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6812_ (.D(_0375_),
    .CLK(net159),
    .Q(\mod.pc_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6813_ (.D(_0376_),
    .CLK(net159),
    .Q(\mod.pc_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6814_ (.D(_0377_),
    .CLK(net153),
    .Q(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6815_ (.D(_0378_),
    .CLK(net152),
    .Q(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6816_ (.D(_0379_),
    .CLK(net153),
    .Q(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0380_),
    .CLK(net195),
    .Q(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0381_),
    .CLK(net195),
    .Q(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0382_),
    .CLK(net194),
    .Q(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0383_),
    .CLK(net194),
    .Q(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0384_),
    .CLK(net194),
    .Q(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0385_),
    .CLK(net179),
    .Q(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0386_),
    .CLK(net180),
    .Q(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0387_),
    .CLK(net179),
    .Q(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0388_),
    .CLK(net178),
    .Q(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0389_),
    .CLK(net178),
    .Q(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0390_),
    .CLK(net177),
    .Q(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0391_),
    .CLK(net177),
    .Q(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6829_ (.D(_0392_),
    .CLK(net172),
    .Q(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6830_ (.D(_0393_),
    .CLK(net173),
    .Q(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6831_ (.D(_0394_),
    .CLK(net173),
    .Q(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6832_ (.D(_0395_),
    .CLK(net172),
    .Q(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6833_ (.D(_0396_),
    .CLK(net172),
    .Q(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6834_ (.D(_0397_),
    .CLK(net172),
    .Q(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6835_ (.D(_0398_),
    .CLK(net173),
    .Q(\mod.instr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6836_ (.D(_0399_),
    .CLK(net177),
    .Q(\mod.instr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6837_ (.D(_0400_),
    .CLK(net177),
    .Q(\mod.instr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6838_ (.D(_0401_),
    .CLK(net187),
    .Q(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6839_ (.D(_0402_),
    .CLK(net164),
    .Q(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6840_ (.D(_0403_),
    .CLK(net165),
    .Q(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6841_ (.D(_0404_),
    .CLK(net164),
    .Q(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6842_ (.D(_0405_),
    .CLK(net192),
    .Q(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6843_ (.D(_0406_),
    .CLK(net192),
    .Q(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6844_ (.D(_0407_),
    .CLK(net192),
    .Q(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6845_ (.D(_0408_),
    .CLK(net194),
    .Q(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6846_ (.D(_0409_),
    .CLK(net175),
    .Q(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6847_ (.D(_0007_),
    .CLK(net170),
    .Q(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6848_ (.D(_0008_),
    .CLK(net175),
    .Q(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6849_ (.D(_0009_),
    .CLK(net168),
    .Q(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6850_ (.D(_0010_),
    .CLK(net168),
    .Q(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6851_ (.D(_0011_),
    .CLK(net170),
    .Q(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6852_ (.D(_0012_),
    .CLK(net168),
    .Q(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6853_ (.D(_0013_),
    .CLK(net169),
    .Q(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6854_ (.D(_0014_),
    .CLK(net171),
    .Q(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6855_ (.D(_0015_),
    .CLK(net169),
    .Q(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6856_ (.D(_0016_),
    .CLK(net168),
    .Q(\mod.instr_2[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6857_ (.D(_0017_),
    .CLK(net170),
    .Q(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6858_ (.D(_0018_),
    .CLK(net175),
    .Q(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6859_ (.D(_0019_),
    .CLK(net170),
    .Q(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6860_ (.D(_0020_),
    .CLK(net183),
    .Q(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6861_ (.D(_0021_),
    .CLK(net163),
    .Q(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6862_ (.D(_0022_),
    .CLK(net183),
    .Q(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6863_ (.D(_0023_),
    .CLK(net165),
    .Q(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6864_ (.D(_0024_),
    .CLK(net164),
    .Q(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6865_ (.D(_0025_),
    .CLK(net164),
    .Q(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6866_ (.D(_0026_),
    .CLK(net165),
    .Q(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6867_ (.D(_0027_),
    .CLK(net152),
    .Q(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6868_ (.D(_0028_),
    .CLK(net151),
    .Q(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6869_ (.D(_0029_),
    .CLK(net151),
    .Q(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6870_ (.D(_0030_),
    .CLK(net151),
    .Q(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6871_ (.D(_0031_),
    .CLK(net151),
    .Q(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6872_ (.D(_0032_),
    .CLK(net163),
    .Q(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6873_ (.D(_0033_),
    .CLK(net163),
    .Q(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6874_ (.D(_0034_),
    .CLK(net188),
    .Q(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6875_ (.D(_0035_),
    .CLK(net187),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6876_ (.D(_0036_),
    .CLK(net152),
    .Q(\mod.ri_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6877_ (.D(_0037_),
    .CLK(net191),
    .Q(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6878_ (.D(_0038_),
    .CLK(net183),
    .Q(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6879_ (.D(_0039_),
    .CLK(net186),
    .Q(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6880_ (.D(_0040_),
    .CLK(net184),
    .Q(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6881_ (.D(_0041_),
    .CLK(net183),
    .Q(\mod.rd_3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6882_ (.D(_0042_),
    .CLK(net193),
    .Q(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6883_ (.D(_0043_),
    .CLK(net176),
    .Q(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6884_ (.D(_0044_),
    .CLK(net176),
    .Q(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6885_ (.D(_0045_),
    .CLK(net175),
    .Q(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6886_ (.D(_0046_),
    .CLK(net166),
    .Q(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6887_ (.D(_0047_),
    .CLK(net167),
    .Q(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6888_ (.D(_0048_),
    .CLK(net166),
    .Q(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6889_ (.D(_0049_),
    .CLK(net166),
    .Q(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6890_ (.D(_0050_),
    .CLK(net166),
    .Q(\mod.ldr_hzd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6891_ (.D(_0051_),
    .CLK(net184),
    .Q(\mod.ldr_hzd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6892_ (.D(_0052_),
    .CLK(net184),
    .Q(\mod.ldr_hzd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6893_ (.D(_0053_),
    .CLK(net185),
    .Q(\mod.ldr_hzd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6894_ (.D(_0054_),
    .CLK(net193),
    .Q(\mod.ldr_hzd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6895_ (.D(_0055_),
    .CLK(net192),
    .Q(\mod.ldr_hzd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6896_ (.D(_0056_),
    .CLK(net190),
    .Q(\mod.ldr_hzd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6897_ (.D(_0057_),
    .CLK(net193),
    .Q(\mod.ldr_hzd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6898_ (.D(_0058_),
    .CLK(net216),
    .Q(\mod.des.des_dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6899_ (.D(_0059_),
    .CLK(net214),
    .Q(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6900_ (.D(_0060_),
    .CLK(net214),
    .Q(\mod.des.des_dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6901_ (.D(_0061_),
    .CLK(net215),
    .Q(\mod.des.des_dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6902_ (.D(_0062_),
    .CLK(net215),
    .Q(\mod.des.des_dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6903_ (.D(_0063_),
    .CLK(net212),
    .Q(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6904_ (.D(_0064_),
    .CLK(net212),
    .Q(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6905_ (.D(_0065_),
    .CLK(net212),
    .Q(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6906_ (.D(_0066_),
    .CLK(net208),
    .Q(\mod.des.des_dout[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6907_ (.D(_0067_),
    .CLK(net209),
    .Q(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6908_ (.D(_0068_),
    .CLK(net212),
    .Q(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6909_ (.D(_0069_),
    .CLK(net209),
    .Q(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6910_ (.D(_0070_),
    .CLK(net213),
    .Q(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6911_ (.D(_0071_),
    .CLK(net122),
    .Q(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6912_ (.D(_0072_),
    .CLK(net122),
    .Q(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6913_ (.D(_0073_),
    .CLK(net114),
    .Q(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6914_ (.D(_0074_),
    .CLK(net112),
    .Q(\mod.registers.r15[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6915_ (.D(_0075_),
    .CLK(net96),
    .Q(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6916_ (.D(_0076_),
    .CLK(net91),
    .Q(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6917_ (.D(_0077_),
    .CLK(net96),
    .Q(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6918_ (.D(_0078_),
    .CLK(net92),
    .Q(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6919_ (.D(_0079_),
    .CLK(net59),
    .Q(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6920_ (.D(_0080_),
    .CLK(net54),
    .Q(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6921_ (.D(_0081_),
    .CLK(net91),
    .Q(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6922_ (.D(_0082_),
    .CLK(net54),
    .Q(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6923_ (.D(_0083_),
    .CLK(net62),
    .Q(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6924_ (.D(_0084_),
    .CLK(net62),
    .Q(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6925_ (.D(_0085_),
    .CLK(net39),
    .Q(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6926_ (.D(_0086_),
    .CLK(net39),
    .Q(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6927_ (.D(_0087_),
    .CLK(net208),
    .Q(\mod.des.des_dout[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6928_ (.D(_0088_),
    .CLK(net208),
    .Q(\mod.des.des_dout[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6929_ (.D(_0089_),
    .CLK(net207),
    .Q(\mod.des.des_dout[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6930_ (.D(_0090_),
    .CLK(net207),
    .Q(\mod.des.des_dout[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6931_ (.D(_0091_),
    .CLK(net210),
    .Q(\mod.des.des_dout[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6932_ (.D(_0092_),
    .CLK(net207),
    .Q(\mod.des.des_dout[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6933_ (.D(_0093_),
    .CLK(net209),
    .Q(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6934_ (.D(_0094_),
    .CLK(net207),
    .Q(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6935_ (.D(_0095_),
    .CLK(net211),
    .Q(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6936_ (.D(_0096_),
    .CLK(net211),
    .Q(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6937_ (.D(_0097_),
    .CLK(net208),
    .Q(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6938_ (.D(_0098_),
    .CLK(net209),
    .Q(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6939_ (.D(_0099_),
    .CLK(net213),
    .Q(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6940_ (.D(_0100_),
    .CLK(net201),
    .Q(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6941_ (.D(_0101_),
    .CLK(net205),
    .Q(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6942_ (.D(_0102_),
    .CLK(net201),
    .Q(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6943_ (.D(_0103_),
    .CLK(net202),
    .Q(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6944_ (.D(_0104_),
    .CLK(net203),
    .Q(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6945_ (.D(_0105_),
    .CLK(net203),
    .Q(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6946_ (.D(_0106_),
    .CLK(net203),
    .Q(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6947_ (.D(_0107_),
    .CLK(net203),
    .Q(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6948_ (.D(_0108_),
    .CLK(net201),
    .Q(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6949_ (.D(_0109_),
    .CLK(net202),
    .Q(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6950_ (.D(_0110_),
    .CLK(net201),
    .Q(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_295 (.ZN(net295));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_296 (.ZN(net296));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_297 (.ZN(net297));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_331 (.ZN(net331));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_332 (.ZN(net332));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_333 (.ZN(net333));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_334 (.ZN(net334));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_335 (.ZN(net335));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_336 (.ZN(net336));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_337 (.ZN(net337));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_338 (.ZN(net338));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_339 (.ZN(net339));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_340 (.ZN(net340));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_341 (.ZN(net341));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_342 (.ZN(net342));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_343 (.ZN(net343));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_344 (.ZN(net344));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_345 (.ZN(net345));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_346 (.ZN(net346));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_347 (.ZN(net347));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_348 (.ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_349 (.ZN(net349));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_350 (.ZN(net350));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_351 (.ZN(net351));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_352 (.ZN(net352));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_353 (.ZN(net353));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_354 (.ZN(net354));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_355 (.ZN(net355));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_356 (.ZN(net356));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_357 (.ZN(net357));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_358 (.ZN(net358));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_359 (.ZN(net359));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_360 (.ZN(net360));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_361 (.ZN(net361));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_362 (.ZN(net362));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_363 (.ZN(net363));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_364 (.ZN(net364));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_365 (.ZN(net365));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_366 (.ZN(net366));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_367 (.ZN(net367));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_368 (.ZN(net368));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_369 (.ZN(net369));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_370 (.ZN(net370));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_371 (.ZN(net371));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_372 (.ZN(net372));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_373 (.ZN(net373));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_374 (.ZN(net374));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_375 (.ZN(net375));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_376 (.ZN(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(io_in[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input12 (.I(io_in[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(io_in[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_in[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(io_in[5]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(io_in[6]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(io_in[7]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(io_in[8]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(io_in[9]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net41),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout41 (.I(net50),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout42 (.I(net45),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net45),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout45 (.I(net49),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net47),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net73),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net55),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net55),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net55),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net61),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net60),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net60),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net60),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net72),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout62 (.I(net65),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net71),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout66 (.I(net70),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net70),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout68 (.I(net70),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net71),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net88),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net77),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net79),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net79),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net87),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout81 (.I(net86),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout82 (.I(net84),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net145),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout90 (.I(net93),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net93),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net99),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net98),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout96 (.I(net98),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout97 (.I(net98),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net109),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net102),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net108),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout103 (.I(net107),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net107),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net107),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net125),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net113),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout114 (.I(net124),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout115 (.I(net119),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout116 (.I(net119),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout117 (.I(net119),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net123),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout120 (.I(net123),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout125 (.I(net144),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net143),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout128 (.I(net143),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net136),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout131 (.I(net135),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net135),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout133 (.I(net135),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout134 (.I(net135),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout135 (.I(net136),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout136 (.I(net142),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout137 (.I(net139),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout138 (.I(net139),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net141),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout143 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net200),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout146 (.I(net147),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net149),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout149 (.I(net162),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout150 (.I(net154),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout151 (.I(net153),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout152 (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout153 (.I(net154),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout154 (.I(net161),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout155 (.I(net156),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net160),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout157 (.I(net160),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout158 (.I(net159),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout159 (.I(net160),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout160 (.I(net161),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout161 (.I(net162),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout162 (.I(net199),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout163 (.I(net199),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout164 (.I(net167),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout165 (.I(net167),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout166 (.I(net167),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout167 (.I(net182),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout168 (.I(net171),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net171),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net171),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout171 (.I(net174),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout172 (.I(net174),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout173 (.I(net174),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout174 (.I(net181),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout175 (.I(net180),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout176 (.I(net180),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout177 (.I(net179),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout178 (.I(net179),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout179 (.I(net180),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout180 (.I(net181),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout181 (.I(net182),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout182 (.I(net198),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout183 (.I(net186),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout184 (.I(net186),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout185 (.I(net186),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout186 (.I(net191),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout187 (.I(net189),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout188 (.I(net189),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout189 (.I(net190),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout190 (.I(net191),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout191 (.I(net197),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout192 (.I(net196),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout193 (.I(net196),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout194 (.I(net196),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout195 (.I(net196),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout196 (.I(net197),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout197 (.I(net198),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout198 (.I(net199),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net200),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout200 (.I(\mod.clk ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout201 (.I(net204),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout202 (.I(net204),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout203 (.I(net205),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(net205),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout205 (.I(net206),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout206 (.I(net218),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout207 (.I(net210),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout208 (.I(net210),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout209 (.I(net210),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout211 (.I(net217),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout212 (.I(net214),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout213 (.I(net214),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net216),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net216),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout216 (.I(net217),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout217 (.I(net218),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout218 (.I(net1),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__RN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__D (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__D (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__D (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__D (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__D (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__D (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__D (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__B1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A3 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A3 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A3 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__B1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__B1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__C (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__C2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__C1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__B1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__B1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__B1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__B1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__B1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__B1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A3 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A3 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__B2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__B1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__I1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__I (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__S (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__S (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I0 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A3 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A3 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A3 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__B (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__B (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__B1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__B2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__S (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__B1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__B2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__B2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A3 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__C (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__I1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__I0 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__C (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__I (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__B1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__B1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__B1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__B1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__B1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__B1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__B1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__B1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__B1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__B1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__B1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__C2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__B1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__B1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__B1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__B1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__B1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__C2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__B1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__B1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__B1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__B1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__B1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__B1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A3 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A3 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__I (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__I1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__B2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__B (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__B1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__B2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__I2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__I3 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__B2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__S (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__S0 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__S0 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__C1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__B1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__C2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__B1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__B1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__B1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__B1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__B1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__B1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__B1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__B1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A4 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A4 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A4 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A4 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__B (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A3 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A4 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A3 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A4 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A3 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A3 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__S (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__S (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__S (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__S (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I0 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__S1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__S1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__S1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__I0 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__B1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__B1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__I1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__I1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A4 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__C (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A3 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__B1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__B1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__B1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__B2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__B (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__I (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__B1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__B1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__B1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__B1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__B1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__B1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I3 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A4 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I3 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__I1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__C2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__B1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__C2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__C1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__B1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__B1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__B1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A3 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__B (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__I1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I0 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A3 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__I0 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A3 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__B (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__B (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A3 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A4 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__B1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I0 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A4 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__B1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__B2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A3 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A4 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__B1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__B2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__B (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I0 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I3 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__S0 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__S0 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__I (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__S0 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__S1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__S1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__B1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__C (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I0 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__B1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__B2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__C (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__I1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__S0 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__S (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__S (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A3 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__I0 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I0 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__I0 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__C1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__B2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__C2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A3 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__C (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I0 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__I (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__B1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__B1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__I (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__B1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__B1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__C1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__B1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__B1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__B1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__C1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__C1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__B1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__C1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__C1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__C1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__B1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__B1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__B1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__B1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__B1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__C2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__C2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__B1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__C2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__B1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__B1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__B1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__B1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__I (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__B1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__B1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__B1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__B1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__B1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__B1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__I (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__B1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__B1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__B1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__B1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__B1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__B (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__B (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__B (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__B1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__C (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__B (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__B (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__C (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A3 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A3 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__B (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__B (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__B (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__B (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A3 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A4 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A3 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__I (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A3 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A4 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__B1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A3 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__B (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__C (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__B1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__B2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__I1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__C (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A3 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A4 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__B1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__B2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A3 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__B2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__B1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__B2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__I2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A3 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__B1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__B2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__B (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__B (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A3 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A3 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A3 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A3 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__B (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A3 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A3 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A4 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__I (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__B (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I3 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__B (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I0 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I0 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__B (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__B (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__B (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__B (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__B2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__S (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__B (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__I (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__B (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I0 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I0 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I0 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A3 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__B (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I3 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__B (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A3 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A3 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__B (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__B1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__B (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__S0 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A3 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A3 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__I (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__S (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__S1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__S1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__B (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__I3 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__S (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I0 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__S0 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__S (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__S (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__I (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A3 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__C (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__B (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I3 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__B2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A3 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A3 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A3 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__B1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__B2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__B2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__B1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__B (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__B2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__C (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__B1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A3 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__B2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A3 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__B (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__C (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__B2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__B (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__B1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__B (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__B2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__C (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__B2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A3 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__I (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__B (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__I0 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__B1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__C (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__B (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__C (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__B (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__C (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__B2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__C (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__S (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A3 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__I (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__B2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__B1 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__B (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A3 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__B2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__C (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__C (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__I (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A3 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__B1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__B1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__B1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__B1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A3 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A4 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__B (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__I0 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__B1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__B (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A3 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A3 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__B1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__C (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A3 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__C (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I0 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I0 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__C (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__C (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__B (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__C (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A3 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__B (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__C (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__C (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__I (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A3 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__C2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__B2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A3 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__C2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A4 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B2 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__B2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__C2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A3 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__B2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A4 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I3 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__B2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A3 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I0 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__C2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A4 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I0 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A4 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__B1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__B1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__C1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__C1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__B1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__B1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__C1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__C1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S0 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__S0 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__S1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__C1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__B1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__B1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__B1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__B1 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__B (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__I (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A3 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__B (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__B1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__I (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__B2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__B (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__B (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__B2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A3 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__B (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__B (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__C (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A3 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__C (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A3 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__C (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A3 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A3 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A3 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__B1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__B (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__B (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__S (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__S (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__B1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__I (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A3 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__B (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__C (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A3 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__B (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__C (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I1 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__B1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__I (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__I1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__C (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__S (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__C (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__I (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__C (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__B1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__I0 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A3 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__B (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__B1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__B1 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__I (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__I (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__I (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__B (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__I (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__I (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A3 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__I (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__B (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__B (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__B (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__I (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__B (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__C (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__B (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__B (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__I (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__I (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A4 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A3 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__B (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__C (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__B (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__B1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__I (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__B1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__I (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__I (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__I (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__I (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__I (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__I (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__I (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__I (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__I (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__I (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__I (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__I (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__I (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__I (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__I (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__I (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__I (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__I (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__I (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__I (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__I (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__I (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__I (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__I (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__I (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__I (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__I (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__I (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__I (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__I (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__I (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__I (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__I (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__B (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__B (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__B (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__I (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__B (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__B (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__B (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__B (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__B (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__B (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__B (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__B (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__I (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__C (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__C (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__C (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__B (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__I (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__I (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__C (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__I (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__B (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__B (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__C (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__B (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__B1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__B (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A3 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A3 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__I (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__B (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I0 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A4 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__I0 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__B (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__B (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__B (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__C (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__C (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__C (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__C (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__I (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__I (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__I (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__I (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__B (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__B (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__B (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A3 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__I (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__I (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__B2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__I (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__B2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__B2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__B2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__I (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B1 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__B2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__B2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__B2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__B2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__I (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__I (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__C (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__C (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__B1 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__I (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__I (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__I (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__B1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__B1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__B1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__B1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__B1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__B1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__I (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__I (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__I (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__B (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__B (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__B (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__B (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__B (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__B (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__B (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__B (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__B (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__B (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__B (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__B (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__B (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__B (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A3 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__I (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__I (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__I (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__B2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__B (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__B (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__B (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__B (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__B2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__B (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__B (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__B (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__B (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__S (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__I (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__S (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__S (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__S (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__S (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__S (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__S (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__S (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__S (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__S (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__S (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__S (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__S (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__I (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__I (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__I (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__I (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__S (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__I (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__S (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__S (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__S (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__S (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__S (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__S (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__S (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__S (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__S (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__S (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__S (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__S (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__I (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__I (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__S (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__S (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__S (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__S (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__S (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__S (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__S (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__S (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__S (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__S (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__S (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__I (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__I (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__B2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__I (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A3 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A3 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__I (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A3 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A3 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__B1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__I (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__C1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__B1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A1 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__I (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A3 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A3 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__I (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A2 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__I (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__I (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__I (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__B1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__B1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__B1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__B1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__C1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__C1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__B1 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__B1 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__C1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__B1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__B1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__B1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__I (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__B1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__I (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__I (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A4 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A4 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__B1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__B1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A2 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__I (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__B1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__B1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__B2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__B2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A3 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__B (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__B (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__C (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B2 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__A1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__I (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__I (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__I (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__I (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__I (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__B (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A3 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__I (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__B (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__I (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__I (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__B (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__B (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__I (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__A2 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__B (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__C (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__I (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__I (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__C (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__B2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__I (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__I (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__B (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__B2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__I (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__I (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A3 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A3 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__I (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A3 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A3 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__B1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__B1 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__B1 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__B1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__B1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__B1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__B1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__B1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A3 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A3 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__B1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__I (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__B1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__B1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__I (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__I (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__B1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__B1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__B1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A3 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A3 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__I (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__I (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__B (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__B (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__I (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A4 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A4 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__I0 (.I(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I0 (.I(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I0 (.I(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__I0 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__I0 (.I(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I0 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__I0 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__I1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I1 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__I1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__I1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__I1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I1 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__I1 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__I1 (.I(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I1 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__I1 (.I(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I1 (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__I0 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I0 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__I (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__B2 (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__B2 (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__I (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__B2 (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__B2 (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__I (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__B2 (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__I (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__B2 (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__B2 (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__B2 (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__I (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__B2 (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__B2 (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__B2 (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__B2 (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A2 (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A2 (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__I (.I(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__I (.I(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A2 (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__C (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__I (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__I (.I(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__I (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I0 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I0 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__I0 (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(\mod.ldr_hzd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(\mod.ldr_hzd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__C2 (.I(\mod.ldr_hzd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(\mod.ldr_hzd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I2 (.I(\mod.ldr_hzd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(\mod.ldr_hzd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I3 (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__B2 (.I(\mod.ldr_hzd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(\mod.ldr_hzd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__I (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__I (.I(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I (.I(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__I (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__I (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__I (.I(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__I (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__I (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__I (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__I (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__I (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__B2 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__A1 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B2 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B2 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__B2 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__B2 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__B2 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__B2 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__B2 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__B2 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__B2 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B2 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B2 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__B2 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__C1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__B2 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__B2 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__B2 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B2 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A3 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__C2 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__B2 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A1 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__B2 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__B2 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__B2 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__B2 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__C2 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A3 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__B2 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__B2 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__B2 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B2 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B2 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A3 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B2 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__C2 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__B2 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B2 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B2 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__B2 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__B2 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B2 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__B2 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A3 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__B2 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__B2 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B2 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__B2 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A3 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B2 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__B2 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__B2 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B2 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__B2 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__B2 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__B2 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__B2 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__B2 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__B2 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__B2 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__B2 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__C1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__B2 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A3 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__B2 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B2 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__B2 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__B2 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__B2 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B2 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__B2 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B2 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__B2 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__B2 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__B2 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__B2 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__B2 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B2 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__B2 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B2 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__B2 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B2 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__B2 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__B2 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__B2 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__B2 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__B2 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B2 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__C1 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__C1 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__B2 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B2 (.I(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__I (.I(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B2 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__B2 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__B2 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__B2 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__B2 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__B2 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__B2 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B2 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__B2 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B2 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A1 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__B2 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__B2 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B2 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__B2 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__B2 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__B2 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__B2 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__B2 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B2 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B2 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A1 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A3 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__C2 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__C1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A3 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__B2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A1 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__B2 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__C2 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__C2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__C1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__B2 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B2 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__B2 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__B2 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__B2 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__B2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__C2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__B2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__B2 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__B2 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B2 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__B2 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__C2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B2 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B2 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__B2 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__B2 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__B2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__B2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__B2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__B2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__B2 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A3 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B2 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__B2 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A3 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__B2 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__B2 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__B2 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__B2 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__B2 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B2 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B2 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__B2 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B2 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B2 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B2 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__B2 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B2 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__B2 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__B2 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B2 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__B2 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__B2 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__C1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__C1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B2 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__I (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B2 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__B2 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__B2 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__C2 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__B2 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__C2 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B2 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__B2 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__B2 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__B2 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__B2 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A3 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__B2 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__B2 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A3 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__B2 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__B2 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B2 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B2 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__B2 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__B2 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__B2 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__B2 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B2 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__B2 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__B2 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A1 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__B2 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__B2 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B2 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__B2 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__B2 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__B2 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__I (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__CLK (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__CLK (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__CLK (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__CLK (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__CLK (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout166_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout170_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout169_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout172_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout173_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__CLK (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout178_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout179_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout176_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout174_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__CLK (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__CLK (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__CLK (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout185_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout189_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout182_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout198_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout199_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout205_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__CLK (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__CLK (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout216_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout206_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1044 ();
 assign io_oeb[0] = net219;
 assign io_oeb[10] = net229;
 assign io_oeb[11] = net230;
 assign io_oeb[12] = net231;
 assign io_oeb[13] = net232;
 assign io_oeb[14] = net233;
 assign io_oeb[15] = net234;
 assign io_oeb[16] = net235;
 assign io_oeb[17] = net236;
 assign io_oeb[18] = net237;
 assign io_oeb[19] = net238;
 assign io_oeb[1] = net220;
 assign io_oeb[20] = net239;
 assign io_oeb[21] = net240;
 assign io_oeb[22] = net241;
 assign io_oeb[23] = net242;
 assign io_oeb[24] = net243;
 assign io_oeb[25] = net244;
 assign io_oeb[26] = net245;
 assign io_oeb[27] = net246;
 assign io_oeb[28] = net247;
 assign io_oeb[29] = net248;
 assign io_oeb[2] = net221;
 assign io_oeb[30] = net249;
 assign io_oeb[31] = net250;
 assign io_oeb[32] = net251;
 assign io_oeb[33] = net252;
 assign io_oeb[34] = net253;
 assign io_oeb[35] = net254;
 assign io_oeb[36] = net255;
 assign io_oeb[37] = net256;
 assign io_oeb[3] = net222;
 assign io_oeb[4] = net223;
 assign io_oeb[5] = net224;
 assign io_oeb[6] = net225;
 assign io_oeb[7] = net226;
 assign io_oeb[8] = net227;
 assign io_oeb[9] = net228;
 assign io_out[0] = net257;
 assign io_out[10] = net267;
 assign io_out[11] = net268;
 assign io_out[12] = net269;
 assign io_out[13] = net270;
 assign io_out[14] = net271;
 assign io_out[15] = net272;
 assign io_out[16] = net273;
 assign io_out[17] = net274;
 assign io_out[18] = net275;
 assign io_out[19] = net276;
 assign io_out[1] = net258;
 assign io_out[2] = net259;
 assign io_out[3] = net260;
 assign io_out[4] = net261;
 assign io_out[5] = net262;
 assign io_out[6] = net263;
 assign io_out[7] = net264;
 assign io_out[8] = net265;
 assign io_out[9] = net266;
 assign la_data_out[0] = net277;
 assign la_data_out[10] = net287;
 assign la_data_out[11] = net288;
 assign la_data_out[12] = net289;
 assign la_data_out[13] = net290;
 assign la_data_out[14] = net291;
 assign la_data_out[15] = net292;
 assign la_data_out[16] = net293;
 assign la_data_out[17] = net294;
 assign la_data_out[18] = net295;
 assign la_data_out[19] = net296;
 assign la_data_out[1] = net278;
 assign la_data_out[20] = net297;
 assign la_data_out[21] = net298;
 assign la_data_out[22] = net299;
 assign la_data_out[23] = net300;
 assign la_data_out[24] = net301;
 assign la_data_out[25] = net302;
 assign la_data_out[26] = net303;
 assign la_data_out[27] = net304;
 assign la_data_out[28] = net305;
 assign la_data_out[29] = net306;
 assign la_data_out[2] = net279;
 assign la_data_out[30] = net307;
 assign la_data_out[31] = net308;
 assign la_data_out[32] = net309;
 assign la_data_out[33] = net310;
 assign la_data_out[34] = net311;
 assign la_data_out[35] = net312;
 assign la_data_out[36] = net313;
 assign la_data_out[37] = net314;
 assign la_data_out[38] = net315;
 assign la_data_out[39] = net316;
 assign la_data_out[3] = net280;
 assign la_data_out[40] = net317;
 assign la_data_out[41] = net318;
 assign la_data_out[42] = net319;
 assign la_data_out[43] = net320;
 assign la_data_out[44] = net321;
 assign la_data_out[45] = net322;
 assign la_data_out[46] = net323;
 assign la_data_out[47] = net324;
 assign la_data_out[48] = net325;
 assign la_data_out[49] = net326;
 assign la_data_out[4] = net281;
 assign la_data_out[50] = net327;
 assign la_data_out[51] = net328;
 assign la_data_out[52] = net329;
 assign la_data_out[53] = net330;
 assign la_data_out[54] = net331;
 assign la_data_out[55] = net332;
 assign la_data_out[56] = net333;
 assign la_data_out[57] = net334;
 assign la_data_out[58] = net335;
 assign la_data_out[59] = net336;
 assign la_data_out[5] = net282;
 assign la_data_out[60] = net337;
 assign la_data_out[61] = net338;
 assign la_data_out[62] = net339;
 assign la_data_out[63] = net340;
 assign la_data_out[6] = net283;
 assign la_data_out[7] = net284;
 assign la_data_out[8] = net285;
 assign la_data_out[9] = net286;
 assign user_irq[0] = net341;
 assign user_irq[1] = net342;
 assign user_irq[2] = net343;
 assign wbs_ack_o = net344;
 assign wbs_dat_o[0] = net345;
 assign wbs_dat_o[10] = net355;
 assign wbs_dat_o[11] = net356;
 assign wbs_dat_o[12] = net357;
 assign wbs_dat_o[13] = net358;
 assign wbs_dat_o[14] = net359;
 assign wbs_dat_o[15] = net360;
 assign wbs_dat_o[16] = net361;
 assign wbs_dat_o[17] = net362;
 assign wbs_dat_o[18] = net363;
 assign wbs_dat_o[19] = net364;
 assign wbs_dat_o[1] = net346;
 assign wbs_dat_o[20] = net365;
 assign wbs_dat_o[21] = net366;
 assign wbs_dat_o[22] = net367;
 assign wbs_dat_o[23] = net368;
 assign wbs_dat_o[24] = net369;
 assign wbs_dat_o[25] = net370;
 assign wbs_dat_o[26] = net371;
 assign wbs_dat_o[27] = net372;
 assign wbs_dat_o[28] = net373;
 assign wbs_dat_o[29] = net374;
 assign wbs_dat_o[2] = net347;
 assign wbs_dat_o[30] = net375;
 assign wbs_dat_o[31] = net376;
 assign wbs_dat_o[3] = net348;
 assign wbs_dat_o[4] = net349;
 assign wbs_dat_o[5] = net350;
 assign wbs_dat_o[6] = net351;
 assign wbs_dat_o[7] = net352;
 assign wbs_dat_o[8] = net353;
 assign wbs_dat_o[9] = net354;
endmodule

