* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5968__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout56_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0074_ net112 mod.registers.r15\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3443__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6845_ _0408_ net194 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6776_ _0339_ net147 mod.pc0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6393__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ mod.registers.r3\[6\] _0979_ _0973_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _2532_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6160__I _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5658_ _2503_ _2500_ _2504_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4156__B1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _0879_ _1581_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5589_ _2107_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5504__I _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3434__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A3 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__A2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3694__I mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4147__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A1 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3673__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _0768_ _1950_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4622__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _3168_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4891_ _1884_ _1874_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3976__A3 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _0196_ net89 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3842_ _0836_ _0837_ _0838_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6375__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _0127_ net78 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4925__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3773_ mod.registers.r6\[5\] _0634_ _0491_ mod.registers.r14\[5\] _0771_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5512_ mod.registers.r6\[2\] _2407_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6492_ _3090_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ mod.registers.r5\[2\] _2350_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4689__B2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ mod.registers.r3\[12\] _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4325_ _1321_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfanout105 net107 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout116 net119 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout127 net143 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout138 net139 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout149 net162 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4256_ _1214_ _1253_ _1195_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4187_ _1181_ _1182_ _1183_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4861__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6155__I mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _0391_ net177 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5169__A2 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4831__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _0325_ net100 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3655__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6065__I mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4065__C1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4514__S _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__A2 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6014__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5409__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3591__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout106_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4135__A3 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__B _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5144__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4110_ _1094_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ mod.pc0\[12\] _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6944__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4041_ _0831_ _0832_ _0833_ _0834_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _2726_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _1929_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4071__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__D _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6348__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4874_ _3189_ _1871_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ _0179_ net110 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3825_ _0819_ _0820_ _0821_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_119_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__I _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _3119_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3756_ _0745_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5571__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ mod.registers.r15\[10\] _3077_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3687_ mod.registers.r6\[2\] _0684_ _0568_ mod.registers.r5\[2\] _0569_ mod.registers.r2\[2\]
+ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_106_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ mod.registers.r4\[15\] _2339_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5323__A2 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5357_ _2176_ _2296_ _2299_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3885__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0459_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _2178_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4239_ _1233_ _1235_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3637__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__B _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__A3 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5562__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__I _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3628__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__C _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4308__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__A1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5139__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _0428_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4590_ _1180_ _1287_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3564__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ mod.registers.r12\[13\] _0504_ _0495_ mod.registers.r15\[13\] _0539_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _2930_ _2939_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3472_ mod.registers.r11\[3\] _3165_ _3167_ mod.registers.r8\[3\] _0470_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _2129_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6191_ _2887_ _2879_ _2889_ _2884_ _2881_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _2057_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3619__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ _0995_ _1017_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_65_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2706_ mod.pc0\[10\] _2710_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4044__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5241__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4926_ mod.pc0\[3\] _1905_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ mod.pc0\[0\] _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ mod.registers.r7\[3\] _0417_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5544__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _1765_ _1785_ _0697_ _0885_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6527_ _3110_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3739_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2358_ _3063_ _3069_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _2320_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6389_ _2932_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4107__I0 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5480__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__A2 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__A1 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__B1 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4274__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5471__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout173_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6253__I _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _2559_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _1706_ _1708_ _1520_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3785__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5691_ mod.registers.r9\[15\] _2521_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4642_ _1130_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4585__I0 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ _1568_ _1569_ _1570_ _0857_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2677_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3524_ mod.registers.r13\[14\] _0490_ _0498_ mod.registers.r4\[14\] _0522_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6243_ _2918_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3455_ _3202_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ mod.des.des_dout\[6\] _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout86_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4657__B _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3386_ _3227_ _3229_ _3236_ _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6239__B1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ _2099_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5056_ _2043_ _0891_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4265__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5462__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4007_ mod.registers.r14\[5\] _3176_ _0710_ mod.registers.r15\[5\] _1005_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__A3 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6163__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _2702_ _2704_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5765__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _1853_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5889_ _2639_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3528__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3528__B2 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6190__A2 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__I _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4591__I3 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__S _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4559__A3 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6685__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6930_ _0090_ net207 mod.des.des_dout\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0021_ net163 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _2517_ _2599_ _2604_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6792_ _0355_ net157 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5747__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ mod.registers.r11\[1\] _2560_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ mod.registers.r9\[10\] _2511_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _1270_ _1620_ _1621_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4183__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4183__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _1142_ _1135_ _0862_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ mod.registers.r6\[15\] _0501_ _0504_ mod.registers.r12\[15\] _0505_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4487_ _1450_ _1473_ _1474_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6226_ _2913_ _2856_ _2914_ _2908_ _2915_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ _3241_ _3229_ _0412_ _3230_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4486__A2 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ mod.des.des_dout\[2\] _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5108_ _2082_ _2092_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _2725_ _2810_ _2813_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5997__I _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4238__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _2024_ _2025_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__B _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3310__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4549__I0 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3980__I mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_223 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_234 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_245 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_256 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_267 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_278 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_289 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3452__A3 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout136_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6154__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _1129_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4165__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ mod.registers.r4\[0\] _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5901__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4986__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _0874_ _1337_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _0482_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4468__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _2741_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3676__B1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__S _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _0073_ net114 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _0407_ net192 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6775_ _0338_ net163 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3987_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5726_ _2530_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5657_ mod.registers.r9\[5\] _2501_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4156__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _1519_ _1593_ _1602_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5588_ _2401_ _2451_ _2456_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3903__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__B2 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _1533_ _1535_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _2674_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3667__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4631__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A4 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4147__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5895__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6300__B _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__B1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__A2 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4890_ _1884_ _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3976__A4 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3841_ mod.registers.r9\[1\] _0423_ _3239_ mod.registers.r10\[1\] _0839_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4490__B _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6375__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _0126_ net74 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3772_ mod.registers.r8\[5\] _3233_ _0632_ mod.registers.r10\[5\] _0770_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5511_ _2353_ _2405_ _2409_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6491_ mod.des.des_dout\[13\] net16 _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6127__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4138__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4689__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _2290_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5605__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _1172_ _1299_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout117 net119 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout128 net143 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout139 net141 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4255_ _1246_ _1251_ _1158_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3649__B1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ mod.registers.r10\[14\] _0895_ _0931_ mod.registers.r9\[14\] _1184_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3416__A3 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__B1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6827_ _0390_ net177 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6366__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6758_ _0324_ net103 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _2499_ _2538_ _2540_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6689_ _0255_ net43 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4129__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5629__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__B1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4065__C2 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5801__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6896__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__B _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3879__B1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ mod.pc_2\[1\] _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5160__I _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__A1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1345_ _1745_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1932_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3803__B1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__A3 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _3190_ _1344_ _1869_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ _0178_ net94 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3824_ mod.registers.r1\[2\] _0747_ _0489_ mod.registers.r13\[2\] _0822_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5020__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3755_ _0746_ _0748_ _0749_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6543_ net8 mod.des.des_dout\[36\] _3106_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _2380_ _3076_ _3079_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3686_ _3154_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5859__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2249_ _2338_ _2342_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4531__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5356_ mod.registers.r3\[5\] _2297_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _1300_ _1301_ _0781_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5287_ _0891_ _2183_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ _1232_ _0963_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ mod.registers.r7\[13\] _0893_ _0918_ mod.registers.r14\[13\] _1166_ _1167_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5070__I mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6036__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5011__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5250__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout216_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ mod.registers.r9\[13\] _0507_ _0513_ mod.registers.r3\[13\] _0538_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3564__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6911__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3471_ mod.registers.r10\[3\] _3161_ _3163_ mod.registers.r9\[3\] _0469_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5155__I _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _1885_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4513__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ mod.des.des_dout\[10\] _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5141_ _2108_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6266__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__B2 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _2058_ _1991_ _1992_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4023_ _0965_ _1019_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3403__I _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__B1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _2714_ _2715_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4044__A3 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4925_ _1896_ _1918_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4234__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4856_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3807_ mod.registers.r5\[3\] _0414_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4787_ _0977_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3555__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ net18 mod.des.des_dout\[28\] _3107_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3738_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6591__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ mod.registers.r15\[3\] _3065_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3669_ _0612_ _0421_ mod.registers.r12\[8\] _0610_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4504__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _2318_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6388_ _1764_ _3017_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5339_ _2108_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6257__A1 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4107__I1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5480__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6771__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__C _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4144__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6934__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3546__A2 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6248__B2 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__I _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout166_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__C _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _1380_ _1707_ _0734_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5690_ _2254_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _1408_ _1410_ _1243_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4734__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _1265_ _1441_ _1443_ _0481_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6311_ _2161_ _2969_ _2972_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3523_ _0500_ _0505_ _0509_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_116_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6487__A1 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3454_ _3223_ _0440_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6242_ _2922_ _2926_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _2855_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3385_ _3230_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6239__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__B2 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _1815_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4229__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ mod.pc_2\[10\] _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ mod.registers.r6\[5\] _0572_ _0716_ mod.registers.r12\[5\] _1004_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5462__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4673__B _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _2703_ _1941_ _2696_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1896_ _1902_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5888_ _2372_ _2647_ _2652_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4839_ mod.ldr_hzd\[13\] _1819_ _1827_ mod.ldr_hzd\[12\] _1822_ mod.ldr_hzd\[15\]
+ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__3528__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ mod.des.des_dout\[21\] net6 _3099_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3308__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6478__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5150__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__C _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5453__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3978__I mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__B _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__I _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _0020_ net183 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5811_ mod.registers.r12\[11\] _2600_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _0354_ net155 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5742_ _2486_ _2558_ _2561_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3758__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _2220_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4707__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4624_ _1477_ _1583_ _1373_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4183__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__A1 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _1268_ _1552_ _1528_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3506_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _1476_ _1480_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4668__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2665_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5132__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _3245_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5343__I _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6156_ _2855_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3368_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _3188_ _1168_ _2091_ _1870_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ mod.pc\[11\] _2766_ _2812_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3299_ _3140_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _2010_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3798__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A2 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5199__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4946__A1 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__B _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4549__I1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5962__B _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5123__A1 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A1 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_224 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_235 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5426__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_246 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_257 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_268 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_279 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5428__I _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4165__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6652__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ _0884_ _0937_ _0943_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _1265_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _2742_ _2743_ _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__B1 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__B2 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6912_ _0072_ net122 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3979__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ _0406_ net192 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _0337_ net190 mod.valid1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ mod.registers.r12\[6\] _0581_ _0583_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6393__A3 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5725_ _2517_ _2544_ _2549_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3600__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__I _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5656_ _2175_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _1354_ _1595_ _1604_ _0869_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5587_ mod.registers.r7\[15\] _2452_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _1340_ _1490_ _1532_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4469_ _1466_ _1218_ _0452_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ mod.instr\[15\] _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3667__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3667__B2 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ mod.pc\[12\] _2679_ _2844_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6081__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4395__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A1 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5647__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3658__B2 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4327__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4083__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4083__B2 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ mod.registers.r7\[1\] _0515_ _0517_ mod.registers.r5\[1\] _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5032__B1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4386__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4630__I0 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ mod.registers.r6\[1\] _2407_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6490_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _2148_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5335__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4138__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5886__A2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5372_ _2288_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4323_ _1300_ _1301_ _1210_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4254_ _0544_ _1170_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4946__B _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__B2 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4310__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ mod.registers.r7\[14\] _0893_ _0929_ mod.registers.r13\[14\] _1183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout61_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4074__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3821__B2 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6698__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _0389_ net178 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5574__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6757_ _0323_ net118 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3969_ mod.registers.r6\[6\] _0684_ _0710_ mod.registers.r15\[6\] _0967_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5708_ mod.registers.r10\[4\] _2539_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6688_ _0254_ net44 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__A1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3316__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6429__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__B2 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6311__B _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout196_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__I _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ mod.pc\[0\] _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _1915_ _1933_ _1916_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3896__I _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3803__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3803__B2 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4872_ _3125_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6611_ _0177_ net110 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4359__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ mod.registers.r7\[2\] _0750_ _0751_ mod.registers.r5\[2\] _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5556__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _3118_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3754_ mod.registers.r7\[7\] _0750_ _0751_ mod.registers.r5\[7\] _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6859__D _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ mod.registers.r15\[9\] _3077_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3685_ _0681_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5859__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ mod.registers.r4\[14\] _2339_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5355_ _2165_ _2296_ _2298_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _0845_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4676__B _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5286_ _2179_ _2052_ _1337_ _2183_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4237_ _1234_ _1018_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4295__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _1163_ _1164_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4099_ mod.registers.r5\[8\] _0897_ _0923_ mod.registers.r2\[8\] _0915_ mod.registers.r11\[8\]
+ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _0372_ net188 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__I _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout111_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout209_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ mod.registers.r6\[3\] _3154_ _3155_ mod.registers.r5\[3\] _3156_ mod.registers.r2\[3\]
+ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _2114_ _2116_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_96_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5171__I _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ mod.funct7\[0\] _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4277__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ _0755_ _0960_ _0962_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4029__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__B2 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _2703_ _2033_ _2707_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4924_ _1752_ _1913_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3806_ _0800_ _0801_ _0802_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4786_ _1773_ _1778_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6736__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _3109_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3737_ _0705_ _0479_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2355_ _3063_ _3068_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3668_ _0612_ _3257_ mod.registers.r11\[8\] _0617_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _2195_ _2326_ _2331_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5701__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _3023_ _3024_ _3022_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3599_ _0444_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6886__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5338_ _2119_ _2257_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _2136_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__B1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__B1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6248__A2 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3482__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout159_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4431__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6759__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4982__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _1355_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _1505_ _1436_ _1508_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4734__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6310_ mod.pc_1\[4\] _2966_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3522_ _0514_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6487__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _3194_ _2924_ _2919_ mod.instr\[2\] _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3453_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4498__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6172_ mod.instr\[6\] _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3384_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5123_ _2098_ _2100_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6239__A2 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__I mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5054_ mod.pc_2\[9\] _2025_ _2027_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5998__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__D _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ mod.registers.r8\[5\] _3168_ _0711_ mod.registers.r9\[5\] _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _2687_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _1896_ _1894_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3776__A3 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5887_ mod.registers.r14\[7\] _2648_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__I _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _1775_ _1826_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4186__B1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ mod.ldr_hzd\[4\] _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6508_ _3088_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6478__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _3057_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4489__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__I _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__B _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4101__B1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5810_ _2515_ _2599_ _2603_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _0353_ net157 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5741_ mod.registers.r11\[0\] _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5672_ _2513_ _2510_ _2514_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4623_ _1389_ _1589_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5904__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3915__B1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4554_ _0882_ _0723_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3505_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4485_ _1109_ _1482_ _0873_ _1395_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5624__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6224_ mod.des.des_dout\[19\] _2866_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout91_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5132__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ _3231_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4340__B1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6155_ mod.instr\[2\] _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ mod.instr_2\[1\] _3218_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4891__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _2083_ _2084_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3298_ mod.registers.r4\[0\] _3144_ _3149_ mod.registers.r1\[0\] _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _2011_ _2015_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4643__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6396__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6396__B2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _2686_ _2689_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput22 net22 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6320__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_225 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_236 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_247 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_258 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_269 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4634__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3988__A3 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__B _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__B _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4270_ _1266_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6947__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3899__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4625__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _0071_ net122 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _0405_ net192 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6378__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ _0336_ net185 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3985_ _0982_ _0445_ mod.registers.r13\[6\] _0583_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ mod.registers.r10\[11\] _2545_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3600__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ _2499_ _2500_ _2502_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _1203_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5586_ _2398_ _2451_ _2455_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4537_ _0732_ _1534_ _0869_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A1 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _0705_ _0844_ _1286_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _2899_ _2891_ _2901_ _2896_ _2893_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3419_ _0411_ _3257_ _3252_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4399_ _3207_ _0859_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4864__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3667__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6185__I mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6069_ _2783_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4616__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3602__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4077__C1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3419__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__B _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__C1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__B _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3512__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4083__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6044__B _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4343__I _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ mod.pc_2\[5\] _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5583__A2 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__I1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ _2353_ _2348_ _2354_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4138__A3 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ _2228_ _2302_ _2307_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5174__I _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4322_ _1290_ _1316_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__A1 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4253_ _1072_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout119 net123 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4184_ mod.registers.r5\[14\] _0898_ _0924_ mod.registers.r2\[14\] _1182_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4074__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__C _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3821__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0388_ net178 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5574__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _0959_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6756_ _0322_ net117 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5707_ _2532_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _0253_ net43 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3899_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _2487_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5569_ _2431_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3888__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4629__S _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__B1 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__B _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6642__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__I _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5014__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3591__A4 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3879__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout189_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4056__A2 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4940_ _1024_ _1914_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__A2 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4871_ _1749_ _1756_ _1855_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _0176_ net110 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ mod.registers.r12\[2\] _0643_ _0644_ mod.registers.r15\[2\] _0820_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ net7 mod.des.des_dout\[35\] _3106_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3753_ _0414_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6472_ _2375_ _3076_ _3078_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3684_ mod.registers.r4\[2\] _0565_ _0566_ mod.registers.r1\[2\] _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _2244_ _2338_ _2341_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3417__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ mod.registers.r3\[4\] _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _1297_ _1299_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _2230_ _2249_ _2250_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4236_ _0766_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4295__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ mod.registers.r13\[13\] _0929_ _0931_ mod.registers.r9\[13\] _1165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4098_ mod.registers.r12\[8\] _0904_ _0917_ mod.registers.r14\[8\] _1096_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4047__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _0371_ net189 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3558__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6739_ _0305_ net116 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6412__B _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__A3 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__I _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4038__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5786__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5538__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__B _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout90 net93 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5717__I _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout104_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5452__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5070_ mod.pc_2\[11\] _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4277__A2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _0767_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__A2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5972_ _2699_ mod.pc0\[9\] _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _1024_ _1914_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4854_ _1757_ _1851_ _1848_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3805_ mod.registers.r4\[3\] _3258_ _3261_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4785_ _1779_ _1780_ _1781_ _1782_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__4201__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3736_ _0723_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6524_ net17 mod.des.des_dout\[27\] _3107_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3960__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ mod.registers.r15\[2\] _3065_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3667_ mod.registers.r6\[8\] _0604_ _0418_ mod.registers.r7\[8\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ mod.registers.r4\[7\] _2327_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6386_ _2933_ _3012_ _3007_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5701__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ mod.instr_2\[4\] _0585_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5337_ _2255_ _2280_ _2285_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5362__I _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5268_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5465__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _0480_ _1027_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _2171_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3476__B1 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3779__B2 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5537__I _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3703__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__B1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6317__B _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3520__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4431__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4195__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _1565_ _1567_ _1379_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4585__I3 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3942__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ mod.registers.r7\[15\] _0516_ _0518_ mod.registers.r5\[15\] _0519_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _2922_ _2925_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _0442_ _3151_ _3186_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6171_ _2873_ _2867_ _2874_ _2872_ _2869_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3383_ mod.instr_2\[11\] _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5122_ mod.rd_3\[2\] _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5447__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _2024_ _2025_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3458__B1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ mod.registers.r4\[5\] _0565_ _0686_ mod.registers.r10\[5\] _1002_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3430__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6703__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _2699_ mod.pc0\[4\] _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4906_ _1897_ _1898_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3630__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3776__A4 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5886_ _2369_ _2647_ _2651_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _1815_ _1830_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4261__I _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4805__S0 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4186__B2 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ mod.ldr_hzd\[5\] _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6507_ _3098_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3719_ mod.registers.r12\[4\] _0716_ _0690_ mod.registers.r14\[4\] _0717_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4699_ _1663_ _1682_ _1696_ _0948_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ mod.des.des_dout\[9\] net7 _3055_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5686__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__I mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6369_ _1780_ _3003_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4436__I _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3340__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5677__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3515__I _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__B2 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout171_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ _2559_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5671_ mod.registers.r9\[9\] _2511_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4622_ _1273_ _1588_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5904__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3915__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4553_ _1546_ _1547_ _1549_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3504_ _0434_ _0435_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4484_ _1413_ _0866_ _1481_ _1397_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5668__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ mod.instr\[19\] _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3435_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3425__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _2860_ _2675_ _2861_ _2859_ _2823_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4340__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4340__B2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3366_ mod.instr_2\[2\] mod.instr_2\[0\] _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _2008_ _2088_ _2089_ _1961_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6085_ _2096_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3297_ _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6093__A1 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _0971_ _1991_ _1992_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5840__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _2688_ _1869_ _0003_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4800__C1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _2638_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3335__I _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4331__B2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__I _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_226 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_237 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_248 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_259 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4634__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6899__CLK net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A2 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5460__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _0070_ net213 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__B1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6841_ _0404_ net164 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__I _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _0002_ _0006_ net218 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3984_ _3173_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5723_ _2515_ _2544_ _2548_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ mod.registers.r9\[4\] _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _1468_ _1219_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5585_ mod.registers.r7\[14\] _2452_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4561__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3364__A2 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _1489_ _1221_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _0845_ _1286_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ mod.des.des_dout\[14\] _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4313__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ mod.registers.r5\[0\] _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4398_ _0875_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _2677_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3349_ mod.instr_2\[2\] mod.instr_2\[0\] _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6068_ _2788_ _2794_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4077__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4077__C2 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3419__A3 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _0982_ _1991_ _1992_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__B1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A3 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__B _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4001__B1 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4304__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4068__B1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A2 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3291__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout134_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6914__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__I _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ mod.registers.r3\[11\] _2303_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4321_ _1317_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _1247_ _1249_ _1090_ _1073_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xfanout109 net125 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4183_ mod.registers.r4\[14\] _0908_ _0926_ mod.registers.r1\[14\] _1181_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6048__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout47_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3282__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _0387_ net179 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5023__A2 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6755_ _0321_ net115 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3967_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _2530_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _0252_ net43 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6594__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3898_ _3155_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5637_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3337__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _2373_ _2439_ _2444_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _1509_ _1510_ _1511_ _1281_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5499_ _2254_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__S0 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__A1 _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__B _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4870_ mod.pc\[0\] _1865_ _1867_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ mod.registers.r9\[2\] _0423_ _0426_ mod.registers.r3\[2\] _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _3117_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3752_ _0417_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6471_ mod.registers.r15\[8\] _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__I mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3683_ mod.registers.r7\[2\] _0679_ _0680_ mod.registers.r3\[2\] _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5422_ mod.registers.r4\[13\] _2339_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4516__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__I1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _2290_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4304_ _1300_ _1234_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5284_ mod.registers.r1\[14\] _2237_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4235_ _1232_ _0963_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3433__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4166_ mod.registers.r11\[13\] _0916_ _0926_ mod.registers.r1\[13\] _1164_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ mod.registers.r7\[8\] _0892_ _0928_ mod.registers.r13\[8\] _1095_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4692__C _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _0370_ net189 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4999_ mod.pc_2\[7\] _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3558__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _0304_ net122 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0235_ net58 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4770__A4 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4507__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5180__A1 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3343__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__B _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5235__A2 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4174__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net93 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4123__B _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4277__A3 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _0993_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _2712_ _2713_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _1915_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _1745_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ mod.registers.r2\[3\] _3250_ _3253_ mod.registers.r11\[3\] _0802_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ mod.ldr_hzd\[0\] _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _3108_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3735_ _0724_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3428__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6454_ _2352_ _3063_ _3067_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3666_ mod.registers.r4\[8\] _3260_ _0621_ mod.registers.r15\[8\] _0664_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5162__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _2188_ _2326_ _2330_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _1765_ _3017_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6632__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ _0447_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5336_ mod.registers.r2\[15\] _2281_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ mod.des.des_dout\[33\] _2207_ _2232_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_102_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5465__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4218_ _1047_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3476__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6782__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _1011_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3476__B2 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ _1143_ _1144_ _1145_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4208__B _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3779__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4728__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3338__I _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3400__A1 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5153__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3703__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3467__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3467__B2 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__I _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4195__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout214_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4788__B _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ _0444_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5463__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ mod.des.des_dout\[5\] _2863_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3382_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5121_ _2099_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6495__S _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _1929_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3458__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3458__B2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5998__A3 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4003_ _0998_ _0999_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6294__I _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5954_ _2700_ _2701_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _1753_ _1899_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3630__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5885_ mod.registers.r14\[6\] _2648_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__B2 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4836_ _1831_ _1832_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__S1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4186__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ mod.ldr_hzd\[6\] _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6506_ mod.des.des_dout\[20\] net5 _3094_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3718_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _1205_ _1254_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ _3056_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5373__I _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3649_ mod.registers.r7\[10\] _0515_ _0517_ mod.registers.r5\[10\] _0647_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6368_ _3005_ _3009_ _3010_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _2262_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6299_ mod.pc_1\[0\] _2679_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3449__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5989__A3 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4110__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3621__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__I _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6678__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5374__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__I _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__B _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout164_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3612__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _2213_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ _3209_ _1611_ _1612_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5365__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3915__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4552_ _1305_ _1302_ _1324_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _3244_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4483_ _1413_ _1433_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3391__A3 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _2911_ _2903_ _2912_ _2908_ _2905_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3434_ _0428_ _0429_ _3245_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_103_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6153_ mod.des.des_dout\[1\] _2856_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _2040_ _2081_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout77_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _2804_ _2806_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ _3145_ _3147_ _3137_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ mod.pc_2\[9\] _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5840__A2 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6820__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5937_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4800__B1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4272__I _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__C2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5868_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ mod.instr_2\[3\] _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5799_ mod.registers.r12\[6\] _2594_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6199__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_227 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_238 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_249 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3351__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4182__I _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5898__A2 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3530__B1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4357__I _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3833__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__B2 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _0403_ net165 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6771_ _0001_ _0005_ net206 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3983_ _0976_ _0977_ _3179_ _0978_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5722_ mod.registers.r10\[10\] _2545_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5653_ _2490_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4604_ _1340_ _1595_ _1598_ _0872_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5584_ _2395_ _2451_ _2454_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _1490_ _1532_ _1354_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4561__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3436__I _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _1460_ _1462_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _2673_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6894__D _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5651__I _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _0482_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3521__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ mod.pc_1\[12\] _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6067_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4077__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3279_ mod.instr_2\[15\] _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4077__B2 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5018_ _1989_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__B2 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4001__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4001__B2 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3760__B1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6057__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6392__I _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__A3 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3291__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5568__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout127_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0631_ _0650_ _1298_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3751__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ _1241_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4182_ _0531_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3282__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _0386_ net180 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ _0320_ net118 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4231__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _0755_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _2497_ _2531_ _2537_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6685_ _0251_ net64 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3897_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5636_ _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5731__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ mod.registers.r7\[7\] _2440_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4518_ _1389_ _1514_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5498_ _2398_ _2391_ _2399_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4449_ _1407_ _1434_ _1446_ _1378_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6531__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4393__S1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6119_ _1957_ _2833_ _2836_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5970__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6522__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A1 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__B _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6202__A2 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3820_ _0814_ _0815_ _0816_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3751_ mod.registers.r9\[7\] _0506_ _0512_ mod.registers.r3\[7\] _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _3064_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ _3138_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5421_ _2236_ _2338_ _2340_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _2288_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _0451_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6297__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__I0 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5283_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ _0755_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4165_ mod.registers.r4\[13\] _0908_ _0895_ mod.registers.r10\[13\] _1163_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4096_ _1092_ _0678_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _0369_ net157 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4204__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ _1752_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _0303_ net46 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5952__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _0944_ _0881_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4755__A2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _0234_ net91 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ _2381_ _2474_ _2477_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5704__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _0165_ net126 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6504__I0 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6904__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4994__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout70 net71 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout81 net86 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout194_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5970_ _2703_ _2021_ _2696_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1897_ _1898_ _1901_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ mod.valid0 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ mod.registers.r6\[3\] _3243_ _3246_ mod.registers.r14\[3\] _0801_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4737__A2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ mod.ldr_hzd\[1\] _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6522_ net16 mod.des.des_dout\[26\] _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3734_ _0728_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4033__C _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ mod.registers.r15\[1\] _3065_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ mod.pc_2\[8\] _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5924__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ mod.registers.r4\[6\] _2327_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _3020_ _3021_ _3022_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3596_ _3202_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5335_ _2249_ _2280_ _2284_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3444__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ _2155_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6111__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4217_ _0965_ _0994_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5197_ _2130_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4673__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3476__A2 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ mod.registers.r10\[12\] _0895_ _0931_ mod.registers.r9\[12\] _1146_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4275__I _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6414__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4079_ mod.registers.r11\[10\] _0577_ _0690_ mod.registers.r14\[10\] _1077_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4425__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__I _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4728__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A1 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3400__A2 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6350__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__A2 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4788__C _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3450_ mod.instr_2\[3\] _0445_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3381_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__B1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _2038_ _1978_ _1981_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3458__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ mod.registers.r2\[5\] _0922_ _3139_ mod.registers.r3\[5\] _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4407__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _2688_ _1923_ _2696_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5080__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4904_ _1038_ _1885_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5884_ _2366_ _2647_ _2650_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3630__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ _1766_ _1820_ _1827_ _1767_ _1823_ _1764_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5383__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ mod.ldr_hzd\[7\] _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3394__A1 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6505_ _3097_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3717_ _3142_ _3170_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _1195_ _1214_ _1253_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ mod.des.des_dout\[8\] net6 _3055_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5135__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3648_ mod.registers.r1\[10\] _0431_ _0433_ mod.registers.r13\[10\] _0646_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6367_ _2666_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3579_ _3165_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5318_ _2260_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6298_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5249_ _2155_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3902__I _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4637__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout157_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4620_ _1355_ _1611_ _1612_ _1615_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4799__B _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6772__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1438_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5474__I _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3502_ _0488_ _0496_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4482_ _1313_ _1365_ _1478_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6314__A1 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ mod.des.des_dout\[18\] _2866_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3433_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6152_ mod.instr\[1\] _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _3192_ _3214_ _3215_ _3198_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_97_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _1209_ _2085_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _2783_ _2808_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3295_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4628__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _1927_ _1448_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4039__B _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5053__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2109_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__B2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4818_ mod.instr_2\[4\] _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5798_ _2503_ _2593_ _2596_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3367__A1 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _1346_ _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6419_ _3046_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput25 net25 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput36 net36 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_228 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_239 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6645__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5559__I _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6241__B1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6795__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3530__B2 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4086__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3833__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5469__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5586__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _0000_ _0004_ net206 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3982_ _0885_ _3180_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _2513_ _2544_ _2547_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _2488_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3349__A1 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__B1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4603_ _1051_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5583_ mod.registers.r7\[13\] _2452_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4534_ _1222_ _1464_ _1469_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4465_ _0735_ _1027_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5932__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ mod.instr\[14\] _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3416_ _0411_ _3242_ _0412_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4396_ _0871_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5510__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3521__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4548__I _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _2064_ _2840_ _2846_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3521__B2 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3347_ mod.instr_2\[1\] _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6668__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2793_ _2030_ _1960_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3278_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5274__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4077__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _1098_ _1099_ _1103_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5577__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ _1851_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _0059_ net214 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4001__A2 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__C _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A3 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3760__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3760__B2 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5063__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4068__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__A1 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3291__A3 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3594__A4 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3537__I _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3751__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3751__B2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6810__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4250_ _1094_ _1107_ _1242_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4368__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4181_ _1177_ _0888_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3282__A3 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ _0385_ net179 mod.instr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6753_ _0319_ net47 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ _0960_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5927__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5704_ mod.registers.r10\[3\] _2533_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6684_ _0250_ net69 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3896_ _0578_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4519__B1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5635_ _2120_ _2458_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3447__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__A3 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5566_ _2370_ _2439_ _2443_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4517_ _1389_ _1442_ _0481_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5497_ mod.registers.r5\[14\] _2392_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5662__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4448_ _1436_ _1437_ _1445_ _1387_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6531__I1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ _1359_ _1365_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ mod.pc_1\[5\] _2834_ _2830_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3910__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6049_ mod.pc\[7\] _2752_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5837__I _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__A2 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3357__I _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6833__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3733__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6522__I1 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__I _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5410__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3750_ mod.registers.r1\[7\] _0747_ _0489_ mod.registers.r13\[7\] _0748_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3681_ _3134_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5420_ mod.registers.r4\[12\] _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _2158_ _2289_ _2295_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__I _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4302_ _3223_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5282_ mod.des.des_dout\[35\] _2178_ _2246_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6513__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ _1215_ _1221_ _1223_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_101_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4164_ mod.registers.r6\[13\] _0903_ _0898_ mod.registers.r5\[13\] _1162_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5229__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _0670_ _0675_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3660__B1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6805_ _0368_ net190 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4997_ _3211_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4204__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5401__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6856__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0302_ net42 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3948_ _0945_ _3214_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6667_ _0233_ net58 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3879_ _0872_ _0873_ _0461_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ mod.registers.r8\[9\] _2475_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5704__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6598_ _0164_ net126 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__B _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5549_ _2430_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__I _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6504__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3651__B1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__I0 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout82 net84 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout93 net99 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__I mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4131__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6729__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout187_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5631__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4434__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6879__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4920_ _1897_ _1898_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4851_ _1759_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5477__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__I _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3802_ mod.registers.r8\[3\] _3232_ _3238_ mod.registers.r10\[3\] _0800_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ mod.ldr_hzd\[2\] _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6521_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3733_ _3194_ _0729_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6452_ _2344_ _3063_ _3066_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5698__A1 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2176_ _2326_ _2329_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3595_ _0564_ _0571_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6383_ _2666_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4370__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__I _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5334_ mod.registers.r2\[14\] _2281_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5940__I _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _1993_ _2185_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4216_ _1155_ _1212_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5196_ _2105_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4147_ mod.registers.r6\[12\] _0903_ _0900_ mod.registers.r3\[12\] _1145_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4078_ mod.registers.r2\[10\] _0569_ _0575_ mod.registers.r9\[10\] _1076_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4425__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5387__I _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__B2 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6719_ _0285_ net48 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5689__A1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3370__I _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3624__B1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5297__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4352__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _3227_ _3229_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6551__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5050_ mod.pc\[10\] _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4104__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__B2 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5852__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4001_ mod.registers.r7\[5\] _3134_ _3148_ mod.registers.r1\[5\] _3166_ mod.registers.r11\[5\]
+ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_78_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4407__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2699_ mod.pc0\[3\] _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4903_ _1038_ _1885_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ mod.registers.r14\[5\] _2648_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _1765_ _1826_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ net14 _1760_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ mod.des.des_dout\[19\] net4 _3094_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3716_ mod.registers.r2\[4\] _0569_ _3144_ mod.registers.r4\[4\] mod.registers.r10\[4\]
+ _0686_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _1420_ _1682_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _3044_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3455__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3647_ mod.registers.r12\[10\] _0643_ _0644_ mod.registers.r15\[10\] _0645_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6332__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _2999_ _3006_ _3008_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ mod.registers.r8\[1\] _0574_ _0575_ mod.registers.r9\[1\] _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_103_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ _2195_ _2268_ _2273_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__I _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _2096_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6096__A1 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ _1950_ _2185_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5843__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _0799_ _2154_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3365__I _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__I _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6087__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4098__B1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6917__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__C _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _1297_ _0676_ _0662_ _0650_ _1298_ _1284_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3501_ mod.registers.r11\[15\] _0497_ _0498_ mod.registers.r4\[15\] _0499_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _0872_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6314__A2 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6220_ mod.instr\[18\] _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4325__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ _0428_ _0429_ _3249_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6151_ _2854_ _2675_ _2857_ _2859_ _2823_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3363_ _3204_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1138_ _2085_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _2788_ _2794_ _2807_ _2805_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3294_ mod.instr_2\[14\] _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5033_ _1873_ _2006_ _2022_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5053__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _2685_ mod.pc0\[0\] _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _2258_ _2583_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6597__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ mod.instr_2\[6\] _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5665__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ mod.registers.r12\[5\] _2594_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3367__A2 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _1213_ _1261_ _1674_ _1212_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6305__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ mod.des.des_dout\[0\] net16 _3045_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ mod.rd_3\[0\] _2852_ _2987_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__S _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5816__A1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_229 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__A2 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__B2 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__B1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4555__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3530__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5807__A1 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__B1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4086__A3 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _3181_ _0580_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5720_ mod.registers.r10\[9\] _2545_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4794__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _2164_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5485__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4546__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _1216_ _1500_ _1599_ _0860_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3349__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__B2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _2390_ _2451_ _2453_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _1520_ _1529_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6299__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A2 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ _2897_ _2891_ _2898_ _2896_ _2893_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3415_ mod.instr_2\[10\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_125_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4395_ _1389_ _1391_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3521__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ mod.pc_1\[11\] _2841_ _2844_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _3195_ _3197_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ mod.pc\[9\] _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__B1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3277_ mod.instr_2\[16\] _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6471__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ _1893_ _1485_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _0058_ net216 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _2375_ _2626_ _2628_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3760__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3751__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _0971_ _0888_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3267__A1 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _0384_ net194 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _0318_ net46 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ _3225_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _2495_ _2531_ _2536_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _0249_ net68 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3895_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__I _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ _2134_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4519__B2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ mod.registers.r7\[6\] _2440_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6635__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ _1290_ _1512_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5164__B _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4447_ _1427_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4378_ _1274_ _1369_ _1372_ _1325_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6785__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _2762_ _2833_ _2835_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3329_ _3131_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _2733_ _2777_ _2778_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4550__S0 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__A3 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3638__I _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3733__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3373__I _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4932__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3421__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout132_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3680_ _0535_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ mod.registers.r3\[3\] _2291_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3724__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5281_ _1179_ _2168_ _2185_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3283__I _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4232_ _1224_ _1225_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ mod.registers.r8\[13\] _0910_ _0920_ mod.registers.r15\[13\] _1161_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5229__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ mod.pc_2\[8\] _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout45_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3660__A1 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3660__B2 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6804_ _0367_ net158 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _1700_ _1703_ _1713_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _0301_ net46 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ _3192_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3412__A1 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0232_ net59 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3878_ _3208_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _2376_ _2474_ _2476_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6597_ _0163_ net139 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5673__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4289__I _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5479_ mod.registers.r5\[10\] _2378_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3921__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__I mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3651__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__B2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout50 net73 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net72 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3706__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4131__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__S _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6431__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3801_ mod.pc_2\[3\] _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5395__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ mod.ldr_hzd\[3\] _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6520_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3732_ mod.funct7\[1\] _3196_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ mod.registers.r15\[0\] _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ mod.pc_2\[9\] _3204_ _0655_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_109_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5698__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ mod.registers.r4\[5\] _2327_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6382_ _2933_ _3006_ _3007_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3594_ _0573_ _0576_ _0579_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _2244_ _2280_ _2283_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4370__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _1138_ _2152_ _2208_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4215_ _1211_ _1171_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3741__I _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _0769_ _2152_ _2168_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ mod.registers.r7\[12\] _0893_ _0926_ mod.registers.r1\[12\] _1144_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A1 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ mod.registers.r6\[10\] _0684_ _0566_ mod.registers.r1\[10\] _0689_ mod.registers.r13\[10\]
+ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5622__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1970_ _1952_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6718_ _0284_ net47 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6499__I _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _0215_ net93 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3916__I _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5310__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5861__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A2 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3624__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3624__B2 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A1 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__B1 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__B1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4104__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6846__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6077__C _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ mod.registers.r5\[5\] _0896_ _3172_ mod.registers.r13\[5\] _0998_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3312__B1 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5852__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5951_ _2698_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4902_ _0961_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5882_ _2361_ _2647_ _2649_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4833_ mod.instr_2\[5\] _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ net15 _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6503_ _3096_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3715_ _0707_ _0708_ _0709_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4695_ _1375_ _1685_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6434_ _3054_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3646_ _0493_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5540__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5951__I _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3577_ _3163_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4995__C _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3551__B1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5316_ mod.registers.r2\[7\] _2269_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2961_ _2962_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6096__A2 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _2127_ _2036_ _2208_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _2131_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4129_ _1022_ _1059_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__I _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5359__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6020__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3646__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__B1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3381__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4098__B2 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5598__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4022__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout212_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _3260_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4480_ _1477_ _1391_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _0413_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5522__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _3212_ _3213_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _2069_ _2072_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1980_ _2048_ _2800_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3293_ mod.instr_2\[15\] _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _1891_ _2007_ _2021_ _1895_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _2676_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5865_ _2400_ _2632_ _2637_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5946__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _1804_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _2499_ _2593_ _2595_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__B _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5761__A1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3466__I _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3772__B1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4678_ _1359_ _1425_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6417_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3629_ _0432_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5513__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5681__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6348_ _2992_ _2996_ _2799_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4297__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ _0445_ _2950_ _2946_ mod.instr\[14\] _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_219 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6241__A2 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4760__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3376__I mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3763__B1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5807__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3818__A1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3818__B2 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout162_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ mod.registers.r7\[6\] _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4243__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _2497_ _2489_ _2498_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _1216_ _0875_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ mod.registers.r7\[12\] _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4532_ _1479_ _1393_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3754__B1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6299__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _1028_ _1031_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6543__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6202_ mod.des.des_dout\[13\] _2888_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3414_ mod.instr_2\[11\] _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4394_ _1317_ _0460_ _1295_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _2038_ _2840_ _2845_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout75_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6064_ _2757_ _2771_ _2782_ _2788_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3276_ mod.instr_2\[17\] _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3809__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__B2 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5015_ _1911_ _1988_ _2004_ _0001_ _2005_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6471__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3285__A2 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6564__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5982__A1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__I _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _0057_ net193 mod.ldr_hzd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ mod.registers.r13\[8\] _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5734__A1 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _2314_ _2457_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3745__B1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3924__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4473__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6214__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6587__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _0383_ net194 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _0317_ net62 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5964__A1 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _0698_ _3191_ _0886_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5496__I _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5702_ mod.registers.r10\[2\] _2533_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6682_ _0248_ net80 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3894_ _3135_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5633_ _2401_ _2480_ _2485_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5564_ _2367_ _2439_ _2442_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5192__A2 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _1266_ _1305_ _1302_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _2248_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__I _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _1439_ _1441_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ mod.pc_1\[4\] _2834_ _2830_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3328_ _3162_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6047_ mod.pc\[6\] _2766_ _2748_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4455__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4550__S1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5955__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _0109_ net202 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3919__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__A4 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A2 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__A2 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4446__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6205__I _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__B1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3421__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout125_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3724__A3 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _0459_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5280_ _2179_ _2093_ _2183_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4231_ _1226_ _1227_ _1057_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4685__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ mod.registers.r12\[13\] _0905_ _0924_ mod.registers.r2\[13\] _0900_ mod.registers.r3\[13\]
+ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_110_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6096__B _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4093_ _1089_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4437__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3660__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6803_ _0366_ net158 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _3126_ _1983_ _1984_ _1986_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__I _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6734_ _0300_ net46 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3946_ _0726_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3412__A2 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _0850_ _0874_ _0854_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6665_ _0231_ net92 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ mod.registers.r8\[8\] _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6596_ _0162_ net138 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6752__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4912__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5547_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _2383_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4429_ _1373_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4428__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout40 net41 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout51 net55 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout62 net65 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout73 net88 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A3 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout95 net98 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4903__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6105__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__B1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4419__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6625__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ _0755_ _0767_ _0781_ _0795_ _0796_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4780_ _1774_ _1775_ _1776_ _1777_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5395__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3731_ _3191_ _0725_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ _0656_ _0657_ _0658_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6344__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _2165_ _2326_ _2328_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6381_ _1766_ _3017_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3593_ _0584_ _0587_ _0588_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ mod.registers.r2\[13\] _2281_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _2140_ _2068_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3705__I0 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4214_ _1211_ _1171_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5194_ _2139_ _1949_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4145_ mod.registers.r4\[12\] _0908_ _0918_ mod.registers.r14\[12\] _1143_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _1072_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5083__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4074__B _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4978_ _0768_ _1950_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6717_ _0283_ net64 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3929_ mod.registers.r2\[15\] _0924_ _0926_ mod.registers.r1\[15\] _0927_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5684__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6335__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6648_ _0214_ net94 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _0145_ net137 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4649__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3932__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6648__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3624__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6798__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3388__B2 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__I _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3560__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3560__B2 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3312__A1 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3312__B2 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout192_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__I _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5950_ _2676_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ mod.pc_2\[2\] _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ mod.registers.r14\[4\] _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4832_ _1824_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3379__A1 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4763_ mod.ins_ldr_3 mod.valid_out3 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ mod.des.des_dout\[18\] net3 _3094_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ mod.registers.r15\[4\] _0710_ _0711_ mod.registers.r9\[4\] mod.registers.r6\[4\]
+ _0684_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4694_ _1395_ _1628_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ mod.des.des_dout\[7\] net5 _3050_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3645_ _0502_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6364_ mod.instr_2\[6\] _2991_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3576_ _3167_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5540__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3551__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _2188_ _2268_ _2272_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3752__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ _1177_ _2957_ _2927_ mod.instr\[20\] _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_114_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ mod.pc_2\[10\] _2198_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3303__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _2126_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _1074_ _1091_ _1110_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4059_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6504__S _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3927__I _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3542__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3542__B2 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4098__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5589__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4270__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4022__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4573__A3 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3430_ _0412_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout205_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3533__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__B _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ mod.funct3\[0\] _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _1177_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3292_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _1882_ _2018_ _2019_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5499__I _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__C _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ _2675_ _2682_ _2684_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ mod.registers.r13\[15\] _2633_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _0613_ _1805_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5210__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ mod.registers.r12\[4\] _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4746_ _0727_ _1741_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5761__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3772__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3772__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _1274_ _1323_ _1325_ _1318_ _1374_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ mod.des.des_counter\[0\] mod.des.des_counter\[1\] mod.des.des_counter\[2\]
+ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3628_ mod.registers.r7\[11\] _0418_ _0415_ mod.registers.r5\[11\] _0626_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5513__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3524__B2 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6347_ mod.ins_ldr_3 _2679_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3559_ mod.registers.r12\[12\] _0504_ _0495_ mod.registers.r15\[12\] _0557_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6278_ _2948_ _2951_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _1914_ _2172_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3288__B1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6033__I _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6836__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3763__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3763__B2 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4488__I _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3392__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5440__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout155_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3567__I _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4600_ _1295_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ _2433_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3754__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4531_ _1380_ _1385_ _1525_ _1526_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3754__B2 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5782__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4462_ _0738_ _1046_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__I1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ mod.instr\[13\] _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4398__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3413_ mod.instr_2\[13\] _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4393_ _1390_ _1027_ _1046_ _1286_ _1271_ _1284_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ mod.pc_1\[10\] _2841_ _2844_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3344_ mod.instr_2\[0\] _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ mod.pc\[9\] _2752_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3275_ _3127_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _0952_ _0957_ _1985_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6709__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout68_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__I0 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3690__B1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6859__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3442__B1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6896_ _0056_ net190 mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _2614_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ _2527_ _2577_ _2582_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _1072_ _1258_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5422__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__I mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3387__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3736__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5489__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4161__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__B1 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _0316_ net62 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _0442_ _0952_ _0957_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ _2493_ _2531_ _2535_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3975__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6681_ _0247_ net102 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3297__I _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3893_ _0885_ _0888_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5632_ mod.registers.r8\[15\] _2481_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ mod.registers.r7\[5\] _2440_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _1232_ _1314_ _1298_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5494_ _2395_ _2391_ _2396_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4445_ _0739_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4152__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__B2 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4376_ _1373_ _1332_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _2826_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3327_ _3170_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2772_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6681__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5687__I _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _0108_ net201 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5955__A2 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _0039_ net186 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4694__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3654__B1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3957__B2 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6422__S _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3709__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ _1226_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5281__B _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _1127_ _1137_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3580__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _0649_ _1084_ _1087_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_370 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _0365_ net154 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _0970_ _0989_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6733_ _0299_ net65 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3412__A3 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _0230_ net96 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3876_ _3213_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _2462_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6595_ _0161_ net138 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6131__I _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4373__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _2286_ _2315_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ _2220_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4125__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4428_ _1283_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4676__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4359_ _1159_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4428__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6029_ mod.pc\[4\] _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4535__B _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__I _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout41 net50 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4600__A2 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net55 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6577__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout96 net98 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4364__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5880__I _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4116__B2 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3627__B1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3661_ mod.registers.r1\[9\] _0510_ _0627_ mod.registers.r13\[9\] _0659_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4355__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ mod.registers.r4\[4\] _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6380_ _3018_ _3019_ _3010_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3592_ mod.registers.r15\[1\] _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _2236_ _2280_ _2282_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _2122_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5855__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3705__I1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4213_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5193_ _2130_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3330__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4075_ _0630_ _1069_ _1071_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5083__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout50_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6126__I _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _1070_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4043__B1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4594__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6716_ _0282_ net68 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3928_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4090__B _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6647_ _0213_ net95 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6335__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3485__I _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6578_ _0144_ net133 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5529_ _2376_ _2418_ _2420_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4649__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__B2 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4821__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3312__A2 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout185_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _1751_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5880_ _2641_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A1 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _1780_ _1826_ _1828_ mod.ldr_hzd\[0\] mod.instr_2\[5\] _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6892__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1750_ _3198_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6501_ _3095_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _3163_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4693_ _1680_ _1396_ _1688_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6317__A2 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4328__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6432_ _3053_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ mod.registers.r9\[10\] _0423_ _0426_ mod.registers.r3\[10\] _0642_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _1820_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3575_ mod.registers.r7\[1\] _3135_ _0572_ mod.registers.r6\[1\] _3139_ mod.registers.r3\[1\]
+ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ mod.registers.r2\[6\] _2269_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3551__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _2940_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ _2197_ _2214_ _2215_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3839__B1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5176_ _2152_ _1913_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4127_ _1111_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5056__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _3222_ _0792_ _0722_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_72_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5695__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6308__A2 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6615__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3542__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5819__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5295__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6765__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4007__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout100_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _3193_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3291_ _3141_ _3130_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_111_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ mod.pc\[8\] _1875_ _1748_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4797__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _2397_ _2632_ _2636_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4814_ _1806_ _1809_ _1810_ _1811_ _0944_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5794_ _2587_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5210__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3772__A2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4676_ _1213_ _1434_ _1259_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6415_ _3042_ _3043_ _2732_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3627_ mod.registers.r9\[11\] _0623_ _0624_ mod.registers.r3\[11\] _0625_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput29 net29 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _0914_ _2851_ _2995_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3558_ mod.registers.r7\[12\] _0516_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _0615_ _2950_ _2946_ mod.instr\[13\] _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6474__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5228_ _2154_ _2006_ _2168_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3288__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3288__B2 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ _2123_ _2135_ _2138_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__B2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4788__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6515__S _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3460__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3763__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6465__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__B _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4453__B _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3848__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout148_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4530_ _1505_ _1527_ _1508_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3754__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6930__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _1452_ _1019_ _1457_ _1458_ _1020_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6200_ _2894_ _2891_ _2895_ _2896_ _2893_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4703__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ _3240_ _3248_ _3256_ _3263_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4392_ _0792_ _0793_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2811_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2725_ _2789_ _2790_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ mod.des.des_counter\[2\] _3121_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _2000_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__I1 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3690__B2 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _2110_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3442__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _0055_ net192 mod.ldr_hzd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3442__B2 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4785__A4 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _2612_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5195__A1 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ mod.registers.r11\[15\] _2578_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4728_ _1670_ _1558_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3745__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _1378_ _1648_ _1650_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3493__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _2043_ _2977_ _2984_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5422__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3736__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__B1 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__A1 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__B2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3220_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3424__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ mod.registers.r10\[1\] _2533_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6680_ _0246_ net105 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3975__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3892_ _0889_ _0887_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ _2398_ _2480_ _2484_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4911__B _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5793__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _2362_ _2439_ _2441_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4513_ _1477_ _1441_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5493_ mod.registers.r5\[13\] _2392_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4444_ _1141_ _1135_ _1132_ _1240_ _0796_ _0600_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4152__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4375_ _0481_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout80_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2824_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3326_ _3142_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4358__B _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _1976_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3663__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6947_ _0107_ net203 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3488__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _0038_ net183 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _2344_ _2613_ _2616_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4143__A2 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5891__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3654__B2 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4715__C _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__B _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3957__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3709__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5118__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6849__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4160_ _1155_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3893__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4091_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_360 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_371 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__B1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _0364_ net162 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _3187_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3944_ _0940_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3948__A2 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6732_ _0298_ net101 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3412__A4 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6663_ _0229_ net91 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3875_ _0847_ _0460_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4641__B _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _2460_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _0160_ net140 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5545_ _2401_ _2424_ _2429_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4373__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3581__B1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5476_ _2381_ _2377_ _2382_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _1303_ _1316_ _1290_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4867__I _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4125__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3333__B1 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _1355_ _0947_ _3209_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ _3159_ _3160_ _3152_ _3153_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _0796_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _1965_ _1966_ _1938_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4061__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout42 net45 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout53 net55 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout75 net77 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3946__I _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout97 net98 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__B1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__I mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5313__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3875__A1 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5616__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__B2 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6433__S _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6232__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3660_ mod.registers.r12\[9\] _0503_ _0621_ mod.registers.r15\[9\] _0658_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3591_ _3128_ _3160_ _3145_ _3174_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5330_ mod.registers.r2\[12\] _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3805__B _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5304__A1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _2197_ _2228_ _2229_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4212_ _1209_ _0464_ _0537_ _0542_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5855__A2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _2160_ _2165_ _2167_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3866__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _1138_ _3223_ _0559_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5607__A2 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4074_ _1069_ _1071_ _0630_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout43_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4043__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__B2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ mod.pc_2\[6\] _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6715_ _0281_ net68 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4594__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _3149_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6142__I _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3858_ _0851_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6646_ _0212_ net89 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5543__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6577_ _0143_ net75 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3789_ mod.registers.r10\[4\] _3239_ _0638_ mod.registers.r4\[4\] _0787_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ mod.registers.r6\[8\] _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _2187_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4282__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__B1 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5534__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4300__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout178_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4830_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5773__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ mod.des.des_dout\[17\] net2 _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3712_ _0589_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3784__B1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4692_ _1193_ _0861_ _1501_ _1689_ _3217_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6431_ mod.des.des_dout\[6\] net4 _3050_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4328__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3643_ _0633_ _0635_ _0637_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5525__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6362_ _1781_ _3003_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _3154_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5313_ _2176_ _2268_ _2271_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6293_ _2955_ _2960_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5828__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__I _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ mod.registers.r1\[9\] _2205_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3839__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3839__B2 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__A2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5175_ _1743_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1121_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6567__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0792_ _0793_ _0722_ _0705_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_72_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4264__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3496__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _1930_ _1935_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _0195_ net113 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4007__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4007__B2 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3766__B1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ _3131_ _3132_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A3 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5931_ _2665_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__A1 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ mod.registers.r13\[14\] _2633_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ mod.ldr_hzd\[4\] _0434_ _1808_ mod.ldr_hzd\[5\] mod.ldr_hzd\[7\] _0424_ _1811_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_5793_ _2585_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4205__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _3194_ _3197_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4675_ _1670_ _1394_ _1499_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _0425_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6414_ _2932_ _3015_ _3036_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ mod.registers.r5\[12\] _0518_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6345_ mod.ri_3 _2852_ _2987_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6276_ _2934_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _3232_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ _0663_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3288__A2 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4808__C _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ mod.registers.r1\[0\] _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109_ _0935_ _1104_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4237__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _1981_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3460__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__B1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__S _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4960__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6330__I _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6732__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4712__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6882__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3451__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__I _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6528__I0 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _1224_ _1225_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4164__B1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3411_ mod.registers.r4\[0\] _3260_ _3262_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4391_ _1282_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _2793_ _2840_ _2843_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3342_ mod.instr_2\[2\] _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ mod.pc\[8\] _2766_ _2748_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3273_ _3126_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5012_ _2001_ _1854_ _2002_ _1961_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3690__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5967__A1 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _2667_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3442__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6894_ _0054_ net193 mod.ldr_hzd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5719__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5845_ _2372_ _2620_ _2625_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _2525_ _2577_ _2581_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6755__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ _1277_ _1724_ _0733_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4942__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6144__A1 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _1653_ _1654_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3609_ _0421_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4589_ _1300_ _0938_ _1301_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ mod.pc_1\[10\] _2982_ _2979_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _1518_ _2935_ _2938_ mod.instr\[7\] _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4458__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__S _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__B1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4697__A1 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4449__B2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6436__S _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3672__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3859__I _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__I _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout160_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ mod.funct7\[2\] _0443_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4621__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3424__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ mod.funct7\[2\] _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ mod.registers.r8\[14\] _2481_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4924__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ mod.registers.r7\[4\] _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4512_ _0863_ _1296_ _1505_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5492_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _1422_ _1272_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4688__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ _1370_ _1240_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3325_ mod.registers.r12\[0\] _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _2750_ _2825_ _2832_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _2742_ _1746_ _1977_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout73_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__A2 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3769__I _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__I mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6946_ _0106_ net203 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _0037_ net191 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ mod.registers.r13\[0\] _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A2 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ _2557_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6117__A1 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__B _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3654__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4603__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3406__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__B _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__I _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4119__B1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3590__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__I _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _1084_ _1087_ _0649_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_350 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_361 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_372 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__B2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _0363_ net155 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _3124_ _1967_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _0297_ net63 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3943_ _0938_ _0936_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _0228_ net96 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6347__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3874_ _0736_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3538__B _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5613_ _2373_ _2468_ _2473_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _0159_ net75 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5309__I _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4213__I _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5544_ mod.registers.r6\[15\] _2425_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3581__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__B2 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5475_ mod.registers.r5\[9\] _2378_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1317_ _1292_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5322__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3333__B2 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4357_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3308_ mod.instr_2\[16\] _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4288_ _1041_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5979__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _2750_ _2752_ _2760_ _2719_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3499__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _0089_ net207 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4061__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout43 net45 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout65 net71 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout76 net77 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4444__S0 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3572__B2 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3875__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5889__I _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__I0 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4461__C _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6816__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _3173_ _0580_ mod.registers.r13\[1\] _0582_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3563__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__I _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ mod.registers.r1\[11\] _2205_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3315__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4211_ mod.pc_2\[13\] _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5191_ mod.registers.r1\[4\] _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3866__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ _0547_ _0550_ _0552_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3330__A4 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073_ _0464_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4815__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4291__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__B1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _1927_ _1635_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5240__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _0280_ net80 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3926_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5791__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6645_ _0211_ net111 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _0852_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ _0142_ net76 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ _0782_ _0783_ _0784_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4878__I _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5527_ _2406_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _2367_ _2363_ _2368_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ _1125_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout200 mod.clk net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout211 net217 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5389_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6256__B1 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3490__B1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5231__A1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6839__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3545__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6508__I _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__S _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__I _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4760_ mod.valid2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3711_ mod.registers.r5\[4\] _0568_ _0574_ mod.registers.r8\[4\] _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3784__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3784__B2 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4691_ _1194_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _3052_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3642_ mod.registers.r4\[10\] _0638_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4328__A3 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3536__A1 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3536__B2 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _3004_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3573_ _0567_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5312_ mod.registers.r2\[5\] _2269_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6292_ mod.funct7\[1\] _2957_ _2927_ mod.instr\[19\] _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5289__A1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3839__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5174_ _2124_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ _0457_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _0965_ _0994_ _1013_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4264__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3472__B1 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5213__A1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5764__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _1931_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _3144_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4972__B1 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4889_ _0830_ _1885_ _1753_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6628_ _0194_ net98 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6559_ _0125_ net74 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__B _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6229__B1 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4007__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3766__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3766__B2 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A4 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5691__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6238__I _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout190_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _2679_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__A2 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _2394_ _2632_ _2635_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3597__I _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ mod.ldr_hzd\[6\] _1807_ _0607_ _0420_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5792_ _2497_ _2586_ _2592_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5746__A2 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3757__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ _1350_ _1737_ _1740_ _3212_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4674_ _1387_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ _1774_ _3034_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3625_ _0422_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6344_ _2961_ _2994_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3556_ mod.registers.r9\[12\] _0507_ _0513_ mod.registers.r3\[12\] _0554_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6275_ _2948_ _2949_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3487_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5226_ _1883_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5682__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5157_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _0457_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ _2068_ _2073_ _2040_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5987__I _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ _0593_ _0598_ _0841_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3996__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3300__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3748__B2 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6537__I1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__I mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3684__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5425__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4306__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4400__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6528__I1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4951__A3 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6557__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6153__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4164__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3410_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout203_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__B2 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1381_ _1386_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__I mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3341_ mod.funct3\[1\] _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _2784_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3272_ _3125_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5664__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ mod.pc0\[7\] _1853_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4219__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ _2667_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ _0053_ net185 mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ mod.registers.r13\[7\] _2621_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5775_ mod.registers.r11\[14\] _2578_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4726_ _1439_ _1268_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3450__I0 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _1427_ _1598_ _1332_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6144__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ mod.registers.r6\[11\] _0604_ _0605_ mod.registers.r14\[11\] _0606_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4588_ _1324_ _1582_ _1584_ _1585_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_1_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4886__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _2981_ _2977_ _2983_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3539_ _0532_ _0533_ _0534_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _2927_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _3200_ _0934_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6189_ _2855_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3666__B1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5407__A1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3969__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__B2 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4570__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A2 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5894__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4449__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__B1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3424__A3 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout153_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5560_ _2433_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4511_ _1505_ _1507_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5491_ _2243_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4442_ _1266_ _1326_ _1321_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4688__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _0863_ _0650_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ mod.pc_1\[3\] _2827_ _2830_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3324_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _2737_ _2773_ _2774_ _2719_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3648__B1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__I _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6062__A1 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6945_ _0105_ net203 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6876_ _0036_ net152 mod.ri_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5827_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__I _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6872__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _2507_ _2565_ _2570_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _1327_ _1546_ _1278_ _1269_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5689_ _2525_ _2520_ _2526_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4679__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5505__I _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__S _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__B1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4064__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3406__A3 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__B1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6071__I _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__C1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4119__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4119__B2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6020__B _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5619__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6745__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__B _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_340 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_351 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_362 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_373 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _1976_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _0296_ net66 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3942_ _0939_ _0937_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6895__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__B1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3819__B _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6661_ _0227_ net111 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ _0851_ _0852_ _0854_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6347__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4358__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ mod.registers.r8\[7\] _2469_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ _0158_ net74 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5543_ _2398_ _2424_ _2428_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3581__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5474_ _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _1422_ _1305_ _1307_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4530__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A2 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _1202_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3307_ _3158_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6026_ _2757_ _2759_ _2751_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5995__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _0088_ net208 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout44 net45 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout55 net61 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6105__B _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6859_ _0019_ net170 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout66 net70 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout77 net79 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout88 net145 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout99 net109 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__S1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3572__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5849__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6768__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__B2 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__I1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3563__A2 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout116_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5145__I _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4512__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _2136_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4141_ _0554_ _0555_ _0556_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5068__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _0420_ _0887_ _0890_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__B2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _1878_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3925_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6713_ _0279_ net117 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6644_ _0210_ net97 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _3193_ _0726_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6575_ _0141_ net75 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ mod.registers.r12\[4\] _0643_ _3247_ mod.registers.r14\[4\] _0785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5526_ _2404_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ mod.registers.r5\[5\] _2364_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5055__I mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _1358_ _1402_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5388_ _2317_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout201 net204 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout212 net214 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4894__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ mod.pc\[2\] _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3490__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3490__B2 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__A1 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3973__I _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3545__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ mod.registers.r3\[4\] _0680_ _0566_ mod.registers.r1\[4\] _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4981__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3784__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _0857_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6933__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3641_ _3261_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3883__I _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3536__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _1782_ _0003_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3572_ mod.registers.r5\[1\] _0568_ _0569_ mod.registers.r2\[1\] _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _2165_ _2268_ _2270_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ _2955_ _2959_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ mod.des.des_dout\[30\] _2207_ _2210_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5173_ _2123_ _2149_ _2150_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _0720_ _0608_ _0887_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4055_ _1036_ _1043_ _1052_ _1032_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3472__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3472__B2 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5213__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4957_ _1086_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3908_ mod.registers.r6\[15\] _0903_ _0905_ mod.registers.r12\[15\] _0906_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4972__A1 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3775__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _0992_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4972__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6627_ _0193_ net110 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3839_ mod.registers.r11\[1\] _0636_ _3247_ mod.registers.r14\[1\] _0837_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6558_ _0124_ net78 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _2345_ _2405_ _2408_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6489_ mod.des.des_counter\[2\] _1872_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6477__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6229__B2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3463__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3766__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4715__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__C1 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout183_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__I0 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A3 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ mod.registers.r13\[13\] _2633_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ mod.ldr_hzd\[10\] _1807_ _1808_ mod.ldr_hzd\[9\] _0424_ mod.ldr_hzd\[11\]
+ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ mod.registers.r12\[3\] _2588_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4403__B1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _1518_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3757__A2 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _1511_ _1669_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6412_ _3040_ _3041_ _2732_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4706__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3624_ mod.registers.r12\[11\] _0503_ _0621_ mod.registers.r15\[11\] _0622_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ net20 _2111_ _2993_ _1346_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3555_ _0547_ _0550_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_115_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ _0607_ _2943_ _2946_ mod.instr\[12\] _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3486_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _2122_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5131__A1 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _2121_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4107_ _0477_ _0609_ _0991_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5087_ _2069_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4038_ _1035_ _0842_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A1 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3996__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1947_ _1948_ _1756_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4945__A1 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3748__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__I _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3684__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__B2 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4936__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__I _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4164__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5361__A1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3340_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3271_ _3123_ _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ mod.pc\[7\] _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3675__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3675__B2 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5416__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3427__A1 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _2667_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6892_ _0052_ net184 mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _2369_ _2620_ _2624_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4927__A1 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ _2523_ _2577_ _2580_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4725_ _1717_ _1718_ _3210_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5328__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__I1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _1439_ _1627_ _1381_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _3246_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4155__A2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1506_ _0827_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6651__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3538_ mod.registers.r4\[13\] _0498_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6326_ mod.pc_1\[9\] _2982_ _2979_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5104__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _2930_ _2937_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3469_ _0465_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _1968_ _2139_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ mod.instr\[10\] _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3666__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3666__B2 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _2118_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3418__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5591__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5894__A2 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__B2 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout146_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5582__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _1383_ _0736_ _0732_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4052__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5490_ _2390_ _2391_ _2393_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4441_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3891__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5885__A2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4372_ _0863_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _2744_ _2825_ _2831_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3323_ _3173_ _3174_ _3170_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ mod.pc\[5\] _2724_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3648__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3648__B2 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout59_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__I _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6944_ _0104_ net203 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4073__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4671__B _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _0035_ net187 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ _2611_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ mod.registers.r11\[7\] _2566_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1270_ _1704_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5688_ mod.registers.r9\[14\] _2521_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4897__I _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _1406_ _1448_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5876__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _2963_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5628__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3639__B2 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4137__I _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3811__B2 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5564__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__B1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3575__C2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4119__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3590__A3 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3878__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_330 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5431__I _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_341 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_352 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_363 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_374 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6044__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _1977_ _1978_ _1979_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _3215_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3802__B2 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__I _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3872_ _0861_ _0864_ _0868_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6660_ _0226_ net97 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _2370_ _2468_ _2472_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4358__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _0157_ net74 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ mod.registers.r6\[14\] _2425_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__A1 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6849__D _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _2213_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _1035_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5858__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ _1127_ _1137_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3306_ mod.instr_2\[17\] _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _0846_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6584__D _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _2740_ _2746_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5341__I _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A2 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _0087_ net208 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6858_ _0018_ net175 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout45 net49 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout56 net60 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__6338__A3 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout67 net70 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout78 net79 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5809_ mod.registers.r12\[10\] _2600_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5546__A1 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6789_ _0352_ net157 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6121__B _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5516__I _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__A2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A2 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3700__S _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout109_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6712__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4512__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3315__A3 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ mod.pc_2\[12\] _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3720__B1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4071_ _1048_ _1064_ _1068_ _0966_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_110_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__I _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6862__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5776__A1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _1759_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3787__B1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _0278_ net117 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3924_ _3156_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5528__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _0209_ net111 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3855_ _0678_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6574_ _0140_ net76 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3786_ mod.registers.r2\[4\] _3251_ _0639_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _2373_ _2412_ _2417_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5456_ _2366_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ _1208_ _0948_ _1403_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5700__A1 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _2318_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout202 net204 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout213 net214 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3711__B1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ _0948_ _1206_ _1257_ _1334_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6256__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ _0826_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__I mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _1744_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3490__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5767__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3778__B1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6735__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6885__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4258__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3481__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5758__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4805__I0 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4981__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _3258_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _3156_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5930__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ mod.registers.r2\[4\] _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6290_ mod.funct7\[0\] _2957_ _2953_ mod.instr\[18\] _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__A2 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _2124_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ mod.registers.r1\[2\] _2137_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4123_ _0564_ _1115_ _1120_ _0966_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_57_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 io_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4054_ _1047_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6608__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3472__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1342_ _1522_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4421__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A2 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _3200_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__I _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _0192_ net112 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3838_ mod.registers.r3\[1\] _0426_ _0644_ mod.registers.r15\[1\] _0836_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4185__B1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _0123_ net85 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3769_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ mod.registers.r6\[0\] _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6488_ _2400_ _3082_ _3087_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6477__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ mod.registers.r5\[1\] _2350_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6229__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3314__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3463__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4412__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3984__I _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3923__C2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3687__C1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3829__I1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout176_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3454__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6900__CLK net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _3236_ _1801_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _2495_ _2586_ _2591_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4403__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _1347_ _1715_ _1735_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3894__I _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6270__I _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _1270_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__B1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6411_ _3026_ _3012_ _3036_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4706__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ _0494_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6342_ _3214_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3554_ _0453_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ _3250_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6273_ _2940_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5614__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _2160_ _2195_ _2196_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _0914_ _1098_ _1099_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5086_ _2070_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4037_ _0599_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4642__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3445__A2 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__C1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6395__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4945__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4939_ _1024_ _1914_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _0175_ net79 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__B _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4633__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3270_ _0000_ mod.des.des_counter\[1\] _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5113__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__I _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3427__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _2666_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _0051_ net184 mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ mod.registers.r13\[6\] _2621_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ mod.registers.r11\[13\] _2578_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4724_ _1638_ _1721_ _0948_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1359_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3606_ _3243_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4586_ _1295_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6325_ _2677_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3537_ _3262_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ mod.instr_2\[6\] _2935_ _2928_ mod.instr\[6\] _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5104__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3468_ mod.registers.r4\[3\] _3143_ _3149_ mod.registers.r1\[3\] _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6946__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _2130_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6187_ _2885_ _2879_ _2886_ _2884_ _2881_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3666__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3399_ _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _1818_ _2100_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3799__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _2055_ _2045_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3418__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5012__C _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5040__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3354__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4606__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4067__C1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5429__I _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6819__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _0739_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4393__I0 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ mod.pc_1\[2\] _2827_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ _3132_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A1 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2770_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3648__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _0103_ net202 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4073__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _0034_ net188 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _2505_ _2565_ _2569_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5573__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _1313_ _1556_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ _2248_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _1486_ _1522_ _1608_ _1635_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5325__A2 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _1324_ _1547_ _1566_ _0847_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6308_ _0799_ _2969_ _2970_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _1750_ _2924_ _2919_ mod.instr\[1\] _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3639__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4836__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6053__A3 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3575__B2 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3590__A4 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_320 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_331 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_342 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_353 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_364 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_375 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3940_ _0724_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6641__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3802__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3871_ _3216_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5004__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5610_ mod.registers.r8\[6\] _2469_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6590_ _0156_ net43 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6791__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _2395_ _2424_ _2427_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5472_ _2376_ _2377_ _2379_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4423_ _1420_ _1412_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3869__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4354_ _1158_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ mod.registers.r6\[0\] _3154_ _3155_ mod.registers.r5\[0\] _3156_ mod.registers.r2\[0\]
+ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ _2753_ _2754_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4294__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _0086_ net39 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _0017_ net170 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout46 net47 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout57 net60 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5808_ _2513_ _2599_ _2602_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout68 net70 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout79 net87 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6788_ _0351_ net146 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3557__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _2556_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3309__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__B1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3761__B _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6363__I _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3796__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3548__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5707__I _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4611__I _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A3 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3720__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__I _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ _1065_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__I _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6273__I _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ _1945_ _1946_ _1963_ _0001_ _1964_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_45_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3787__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ _0277_ net105 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3923_ mod.registers.r11\[15\] _0916_ _0918_ mod.registers.r14\[15\] mod.registers.r15\[15\]
+ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__3787__B2 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6642_ _0208_ net111 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3854_ mod.funct3\[0\] _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3539__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3846__B _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _0139_ net82 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3785_ mod.registers.r9\[4\] _0506_ _0636_ mod.registers.r11\[4\] _0783_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ mod.registers.r6\[7\] _2413_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5455_ _2175_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _1352_ _1246_ _1251_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5700__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout203 net205 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout214 net216 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3711__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _1200_ _1201_ _3210_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3711__B2 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__I _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4268_ _1035_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6500__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ mod.valid2 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__B1 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4019__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6183__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3778__A1 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6909_ _0069_ net209 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__B2 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5527__I _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5262__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4258__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3481__A3 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3510__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__I1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5437__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ _3155_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3941__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ _1122_ _2181_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _1116_ _1117_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5105__C _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _1048_ _0698_ _1049_ _1050_ _0824_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__I _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 io_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _1878_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3906_ _0715_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4886_ _1861_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _0191_ net40 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3837_ _0831_ _0832_ _0833_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4185__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4185__B2 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _0122_ net82 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3768_ mod.pc_2\[6\] _0594_ _0760_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5507_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ mod.registers.r15\[15\] _3083_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3699_ _3180_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__B _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _2221_ _2302_ _2306_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3696__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__C _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6127__B _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6702__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4870__B _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A3 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4176__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6852__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3505__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__B1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__C2 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3439__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__B _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__A3 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout169_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _0851_ _1336_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _1370_ _1283_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4167__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _1775_ _3034_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4167__B2 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3622_ _0603_ _0606_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5903__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3553_ mod.registers.r4\[12\] _0498_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6272_ _2941_ _2947_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3484_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ mod.registers.r1\[7\] _2166_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3415__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ mod.des.des_dout\[21\] _2125_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__D _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4105_ _1100_ _1101_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_96_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5085_ _2055_ _2045_ _2060_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6092__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ _1023_ _1032_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6725__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__C2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _2723_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _1930_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5077__I mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _0174_ net79 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ net6 mod.des.des_dout\[34\] _3106_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__B1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4330__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6083__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5830__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4633__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__B1 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6320__B _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5450__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6890_ _0050_ net166 mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _2366_ _2620_ _2623_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6281__I _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _2519_ _2577_ _2579_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _1245_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6129__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _1285_ _1372_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5888__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3605_ mod.registers.r8\[11\] _3234_ _0602_ mod.registers.r10\[11\] _0603_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4585_ _1232_ _0767_ _1240_ _1314_ _0826_ _0846_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5625__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2024_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4560__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3536_ mod.registers.r2\[13\] _0485_ _0497_ mod.registers.r11\[13\] _0534_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6255_ _2930_ _2936_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ mod.registers.r7\[3\] _3135_ _3138_ mod.registers.r3\[3\] _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4312__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _2179_ _1967_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6186_ mod.des.des_dout\[9\] _2876_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3398_ _3235_ _3230_ _3249_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ mod.rd_3\[0\] _2101_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ mod.pc_2\[10\] _0891_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _1014_ _1015_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__B1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4000__B1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__C _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__B1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4067__C2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3939__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4790__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6050__B _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout201_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _1366_ _0631_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4393__I1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6570__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3321_ _3152_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _2756_ _2771_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6276__I _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _0102_ net201 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _0033_ net163 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5824_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ mod.registers.r11\[6\] _2566_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4706_ _1296_ _1548_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5686_ _2523_ _2520_ _2524_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6913__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _1609_ _1618_ _1619_ _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4128__A4 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _0842_ _0825_ _0459_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6307_ mod.pc_1\[3\] _2966_ _2964_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3519_ _0414_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1284_ _1282_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5089__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _2670_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ mod.instr\[5\] _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5261__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__A2 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6277__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_310 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3513__I _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_321 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_332 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_343 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_354 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_365 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_376 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout151_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _0866_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5004__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6936__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4212__B1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ mod.registers.r6\[13\] _2425_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4763__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ mod.registers.r5\[8\] _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3971__C1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__I _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4422_ _1341_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4515__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A3 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4353_ _3212_ _1338_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6268__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3304_ _3152_ _3153_ _3137_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6268__B2 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _0701_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout64_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6925_ _0085_ net39 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6856_ _0016_ net168 mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net60 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5807_ mod.registers.r12\[9\] _2600_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6787_ _0350_ net149 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3999_ mod.pc_2\[5\] _0594_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3557__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5738_ _2557_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4203__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _2509_ _2510_ _2512_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4506__B2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3714__C1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6259__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6259__B2 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3508__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A1 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3720__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _3124_ _1949_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6710_ _0276_ net106 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3922_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3787__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6641_ _0207_ net40 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3539__A2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6572_ _0138_ net128 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3784_ mod.registers.r5\[4\] _0751_ _0644_ mod.registers.r15\[4\] _0782_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ _2370_ _2412_ _2416_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4023__B _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5454_ _2362_ _2363_ _2365_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _1246_ _1251_ _1352_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5385_ _2315_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4336_ _0942_ _1258_ _1263_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3711__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout204 net205 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout215 net216 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4249__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4267_ _0828_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6006_ _1965_ _1966_ _1904_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4198_ _0544_ _1171_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3475__B2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5216__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _0068_ net212 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3778__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _0402_ net164 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4188__C1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3702__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6374__I _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6404__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__I2 mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6323__B _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4718__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout114_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__A2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ mod.des.des_dout\[23\] _2125_ _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4121_ mod.registers.r12\[9\] _0904_ _0919_ mod.registers.r15\[9\] _1119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _0725_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3457__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6284__I _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _1758_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3905_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _1866_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4709__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _0190_ net38 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ mod.registers.r4\[1\] _0638_ _0639_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _0121_ net85 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3767_ _0761_ _0762_ _0763_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5506_ _2403_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6486_ _2397_ _3082_ _3086_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3698_ _0443_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _2143_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5363__I _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5368_ mod.registers.r3\[10\] _2303_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3696__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3696__B2 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4319_ _0797_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3448__A1 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3620__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5982__B _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4176__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3687__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3687__B2 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3722__S _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__B2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _0884_ _1546_ _1384_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3621_ _3203_ _0611_ _0614_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4167__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ _0548_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6340_ _0851_ _1760_ _2668_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ _1802_ _2943_ _2946_ mod.instr\[11\] _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3483_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3678__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3678__B2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5153_ _3224_ _2127_ _2128_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__I _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ mod.registers.r1\[8\] _0925_ _0919_ mod.registers.r15\[8\] _1102_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5084_ _2057_ _2059_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _0480_ _0811_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6092__A2 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3850__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1747_ _1864_ _2109_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ mod.pc_2\[4\] _1122_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _1747_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6607_ _0173_ net77 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5355__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ mod.registers.r4\[2\] _3259_ _0639_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _1772_ _1789_ _0971_ _0476_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _3116_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _3062_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3606__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4330__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__B _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3841__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3841__B2 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4397__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5268__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4321__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout181_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4347__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ mod.registers.r13\[5\] _2621_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5585__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ mod.registers.r11\[12\] _2578_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _1091_ _1643_ _1089_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _1285_ _1361_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5888__A2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3604_ _3238_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _0795_ _1366_ _1363_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6323_ _1092_ _2977_ _2980_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3535_ mod.registers.r6\[13\] _0501_ _0492_ mod.registers.r14\[13\] _0533_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3426__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _2933_ _2935_ _2928_ mod.instr\[5\] _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3466_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1883_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ mod.instr\[9\] _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3397_ _3241_ _3228_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5136_ _1821_ _2100_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _2008_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4076__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6842__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _0781_ _1012_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5812__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3823__B2 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5969_ _2699_ mod.pc0\[8\] _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__B2 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__A3 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3336__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4839__B1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3511__B1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A4 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4067__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4067__B2 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3578__B1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__B _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4790__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5726__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6715__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__I2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3320_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3750__B1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__S _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__A1 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _0101_ net205 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6872_ _0032_ net163 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ _2120_ _2583_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5558__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3569__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _2503_ _2565_ _2568_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4230__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ _1663_ _1702_ _1609_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5685_ mod.registers.r9\[13\] _2521_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1624_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4533__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5730__A1 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _1422_ _1512_ _1513_ _1312_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6306_ _2848_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3518_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4696__B _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _1207_ _1492_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _2922_ _2923_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3449_ mod.funct3\[2\] _0446_ _3201_ mod.instr_2\[1\] _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _2870_ _2867_ _2871_ _2872_ _2869_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ mod.ins_ldr_3 mod.valid_out3 net15 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4049__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6099_ _2683_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__A1 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6210__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6738__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3775__B _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6888__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6377__I _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6277__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_300 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_311 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_322 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_333 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_344 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5088__I0 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_355 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_366 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6326__B _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4212__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4212__B2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6061__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__I _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3971__B1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5470_ _2349_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3971__C2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _1205_ _1412_ _1415_ _1417_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4515__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4352_ _0865_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3303_ _3128_ _3129_ _3131_ _3146_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6287__I _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4283_ _0737_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3704__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _2740_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout57_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _0084_ net62 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6855_ _0015_ net169 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ _2509_ _2599_ _2601_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout59 net60 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4203__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _0349_ net147 mod.pc0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3998_ _0774_ _0779_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5737_ _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ mod.registers.r9\[8\] _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5703__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _1204_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4506__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5599_ _2353_ _2461_ _2465_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3714__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3714__C2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__I mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6259__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6560__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5942__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__B1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5170__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3800__S0 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__S _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6056__B _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6903__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1956_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _0589_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _0206_ net40 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3852_ _3191_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ _0137_ net86 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5933__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5522_ mod.registers.r6\[6\] _2413_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6489__A2 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5453_ mod.registers.r5\[4\] _2364_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5914__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _1377_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5384_ _2114_ _2116_ _2118_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4335_ _1264_ _1280_ _1331_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout205 net206 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout216 net217 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _0856_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4121__B1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _1193_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__A2 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6907_ _0067_ net209 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__I _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _0401_ net187 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4188__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4188__C2 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _0335_ net48 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3609__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A3 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__I mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__I3 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3519__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6340__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ mod.registers.r6\[9\] _0902_ _0909_ mod.registers.r8\[9\] _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4794__B _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4051_ _0683_ _0695_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_96_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _1001_ _1002_ _1006_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _0572_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4884_ mod.pc0\[1\] _1876_ _1877_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6623_ _0189_ net51 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5906__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4709__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3835_ mod.registers.r2\[1\] _3251_ _0431_ mod.registers.r1\[1\] _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _0120_ net82 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3766_ mod.registers.r7\[6\] _0515_ _0517_ mod.registers.r5\[6\] _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3393__A1 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5505_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ mod.registers.r15\[14\] _3083_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ _0685_ _0687_ _0688_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _2345_ _2348_ _2351_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5367_ _2214_ _2302_ _2305_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4893__A1 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3696__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ _1306_ _0662_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5298_ _2259_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ _1089_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4645__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3448__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__B2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3620__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3339__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3908__B1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3687__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4884__B2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6334__B _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _0615_ _0616_ mod.registers.r11\[11\] _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3551_ mod.registers.r6\[12\] _0501_ _0492_ mod.registers.r14\[12\] _0549_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5464__I _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6313__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _2918_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3482_ _0464_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ mod.des.des_dout\[28\] _2151_ _2191_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3678__A2 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5152_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ mod.registers.r6\[8\] _0902_ _0894_ mod.registers.r10\[8\] _1101_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ mod.pc_2\[12\] _1177_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3712__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4034_ _1029_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _2721_ _2722_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5639__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ mod.pc_2\[4\] _1122_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6606_ _0172_ net77 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3818_ mod.registers.r2\[2\] _0483_ _0636_ mod.registers.r11\[2\] _0816_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4798_ _1779_ _1787_ _1785_ _1780_ _1788_ _1781_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__3366__A1 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6771__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6537_ net5 mod.des.des_dout\[33\] _3112_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3749_ _0430_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _2372_ _3070_ _3075_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _2320_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6399_ _2684_ _3032_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3669__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4330__A3 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5043__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__A1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout174_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _2559_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5585__A2 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _1663_ _1717_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6794__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _1238_ _1258_ _1630_ _1090_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3603_ _0521_ _0531_ _0544_ _0561_ _0563_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4583_ _1571_ _1578_ _1580_ _3217_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3707__I _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ mod.pc_1\[8\] _2973_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3534_ mod.registers.r8\[13\] _0487_ _0508_ mod.registers.r10\[13\] _0532_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3465_ _3221_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5922__I _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _2129_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6184_ _2882_ _2879_ _2883_ _2884_ _2881_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ mod.registers.r6\[0\] _3244_ _3247_ mod.registers.r14\[0\] _3248_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ mod.rd_3\[1\] _2101_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _2052_ _1734_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5273__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__I0 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _0794_ _0723_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _2705_ _2004_ _2711_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5576__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _1105_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5899_ _2639_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3511__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3511__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3352__I _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6667__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3578__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3578__B2 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4393__I3 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3750__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3750__B2 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__I0 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _0100_ net201 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ _0031_ net151 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4307__B _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5189__I _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5822_ _2527_ _2605_ _2610_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3569__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5753_ mod.registers.r11\[5\] _2566_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3569__B2 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5917__I _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _1452_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _2243_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _1479_ _1628_ _1631_ _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1264_ _1560_ _1563_ _1418_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _0813_ _2849_ _2968_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _0417_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4497_ _1454_ _1493_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5652__I _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6236_ _3196_ _2671_ _2919_ mod.instr\[0\] _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3448_ mod.instr_2\[2\] mod.instr_2\[0\] _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5494__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4268__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _2858_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ mod.instr_2\[11\] _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _1831_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6098_ _2819_ _2820_ _2751_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4049__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ mod.pc0\[10\] _1958_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3900__I _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__I _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4221__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__C _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3347__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4178__I _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_301 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_312 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_323 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_334 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_345 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_356 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_367 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5788__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4460__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4212__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout137_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _0869_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4515__A3 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__B _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _1347_ _1348_ _1338_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3302_ _3128_ _3130_ _3152_ _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _0733_ _1269_ _1275_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4279__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _2741_ _2745_ _2753_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_98_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6923_ _0083_ net62 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4451__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _0014_ net171 mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout38 net41 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ mod.registers.r12\[8\] _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6785_ _0348_ net150 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4203__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _0965_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _2286_ _2458_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5667_ _2490_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4618_ _1610_ _1614_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5703__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ mod.registers.r8\[1\] _2463_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3714__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3714__B2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _0795_ _0812_ _0862_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5382__I _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6219_ _2909_ _2903_ _2910_ _2908_ _2905_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4514__I0 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6705__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3786__B _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__S1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5458__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6337__B _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4984__A3 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3851_ _0737_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6072__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5467__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _0136_ net80 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3782_ _0769_ _0678_ _0774_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _2367_ _2412_ _2415_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _2349_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4403_ _1378_ _1388_ _1393_ _1395_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5383_ _2314_ _2107_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4334_ _0945_ _0855_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout206 net218 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout217 net218 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4265_ _0940_ _1259_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4121__A1 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _2726_ _2728_ _1880_ _2734_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4121__B2 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ _0525_ _0530_ _1176_ _1191_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6728__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3475__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ _0066_ net208 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6878__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _0400_ net177 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__S0 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__B2 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6768_ _0334_ net47 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3935__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _2509_ _2544_ _2546_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6699_ _0265_ net66 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3625__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5860__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4456__I _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3360__I _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5996__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6340__A2 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4103__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ _0564_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4103__B2 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3457__A3 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5603__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ _0000_ mod.des.des_counter\[1\] _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__C1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3903_ mod.registers.r5\[15\] _0898_ _0900_ mod.registers.r3\[15\] _0901_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4883_ _1759_ _1878_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _0188_ net51 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3834_ mod.registers.r6\[1\] _3244_ _0643_ mod.registers.r12\[1\] _0832_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5906__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _0119_ net133 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3765_ mod.registers.r9\[6\] _0623_ _0624_ mod.registers.r3\[6\] _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4969__C _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4590__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6484_ _2394_ _3082_ _3085_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3696_ mod.registers.r13\[2\] _0689_ _0690_ mod.registers.r14\[2\] _0693_ _0694_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ mod.registers.r5\[0\] _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5366_ mod.registers.r3\[9\] _2303_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6550__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _1306_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _1231_ _1237_ _1244_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4276__I _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4179_ _0889_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__B1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3620__A3 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3908__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3908__B2 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__B _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5570__I _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__B1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A3 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout217_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3550_ mod.registers.r8\[12\] _0487_ _0508_ mod.registers.r10\[12\] _0548_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3481_ _0442_ _0467_ _0475_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_6_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _2171_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5151_ _2129_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ mod.registers.r3\[8\] _0899_ _0909_ mod.registers.r8\[8\] _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5082_ _2052_ _1406_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _0706_ _0477_ _1030_ _3199_ _0811_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2703_ _2091_ _2707_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4935_ _1884_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _1850_ _1856_ _1863_ _1847_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6605_ _0171_ net83 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6916__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3817_ mod.registers.r6\[2\] _0634_ _0491_ mod.registers.r14\[2\] _0815_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _1782_ _1789_ _0973_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4699__C _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3366__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ mod.registers.r12\[7\] _0502_ _0494_ mod.registers.r15\[7\] _0746_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6536_ _3115_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _0631_ _0650_ _0662_ _0676_ _0563_ _0600_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6467_ mod.registers.r15\[7\] _3071_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _2318_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6398_ _1770_ _3028_ _3029_ _3012_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3669__A3 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5349_ _2149_ _2289_ _2294_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4079__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5815__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__B1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6154__C _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6240__A1 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4554__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4609__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3817__B1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__B _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout167_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4720_ _1245_ _1133_ _1716_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _1089_ _1501_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3602_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4545__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _1573_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3533_ _0525_ _0530_ _3205_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6321_ _2963_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _2669_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3464_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _2160_ _2176_ _2177_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4819__I mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _2858_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3395_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _1927_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4320__I1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__B2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ _2706_ mod.pc0\[7\] _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ _3211_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5898_ _2386_ _2653_ _2658_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4849_ _1763_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ mod.des.des_counter\[2\] _1945_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3633__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3511__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6461__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4775__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3578__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4527__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3750__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3502__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4550__I1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4058__A3 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _0030_ net151 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ mod.registers.r12\[15\] _2606_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3569__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _2499_ _2565_ _2567_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _1235_ _1616_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4323__B _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _2519_ _2520_ _2522_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3718__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _1234_ _1018_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5191__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _1541_ _1562_ _1203_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6304_ mod.pc_1\[2\] _2966_ _2964_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3516_ mod.registers.r1\[15\] _0511_ _0513_ mod.registers.r3\[15\] _0514_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4496_ _1454_ _1493_ _1204_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__B _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _2915_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3447_ _3174_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3453__I _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ mod.des.des_dout\[4\] _2863_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3378_ mod.instr_2\[10\] _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _2097_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6097_ _2819_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4049__A3 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5048_ _1893_ _1659_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input12_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4284__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3829__S _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3732__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3363__I _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6784__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_302 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_313 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_324 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_335 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_346 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_357 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_368 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4599__I1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__A2 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5173__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ _3193_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3723__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ _3132_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3273__I _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _1345_ _2743_ _2750_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6922_ _0082_ net54 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4451__A3 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _0013_ net169 mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5804_ _2587_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _0347_ net148 mod.pc0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _0766_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5735_ _2527_ _2550_ _2555_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3411__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6657__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3962__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _2488_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4617_ _1610_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5597_ _2345_ _2461_ _2464_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4911__A1 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3714__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1506_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4479_ _0739_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ mod.des.des_dout\[17\] _2900_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4514__I1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _1856_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3911__I _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4442__A3 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__I _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__A2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4115__C1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3469__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__A1 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ _0739_ _0798_ _0827_ _0829_ _0843_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ _0775_ _0776_ _0777_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ mod.registers.r6\[5\] _2413_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3944__A2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _2347_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4402_ _1352_ _1396_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5382_ _2103_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4333_ _1281_ _1311_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout207 net210 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__6497__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout218 net1 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4264_ _0941_ _1261_ _0947_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6003_ _2733_ _2736_ _2738_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4121__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _1176_ _1179_ _1180_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout62_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _0065_ net212 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3632__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3632__B2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6836_ _0399_ net177 mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__S1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _0333_ net64 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ _0585_ _0586_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3396__B1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3935__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5718_ mod.registers.r10\[8\] _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6698_ _0264_ net66 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5649_ mod.registers.r9\[3\] _2491_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3906__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4112__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3641__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5996__C _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__CLK net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__A1 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5128__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4351__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6348__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__A1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4103__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout197_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__A2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5064__B1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5603__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4951_ _1942_ _1943_ _1944_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4382__I _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__C2 mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3902_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4882_ mod.pc\[1\] _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6621_ _0187_ net58 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ mod.registers.r8\[1\] _0486_ _0433_ mod.registers.r13\[1\] _0831_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6552_ _0118_ net141 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3764_ mod.registers.r1\[6\] _0431_ _0627_ mod.registers.r13\[6\] _0762_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _2258_ _2315_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5119__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ mod.registers.r15\[13\] _3083_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3695_ _0691_ _3178_ _3179_ _3182_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6102__I _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5365_ _2204_ _2302_ _2304_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3550__B1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4316_ _1094_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4247_ _1074_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6845__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _3205_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3605__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5388__I _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4292__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6819_ _0382_ net194 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3908__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4030__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3636__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5530__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__B1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__I _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__B2 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5833__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5597__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6010__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4021__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__B1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3480_ _0444_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4324__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6868__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _1750_ _3201_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ mod.registers.r4\[8\] _0907_ _0930_ mod.registers.r9\[8\] _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5081_ _1872_ _2053_ _2066_ _3126_ _2067_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4088__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ _0467_ _0475_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_96_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3835__B2 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ mod.pc0\[13\] _2685_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _1927_ _1538_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _1758_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5936__I _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6604_ _0170_ net126 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3816_ mod.registers.r8\[2\] _3233_ _0632_ mod.registers.r10\[2\] _0814_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4012__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1792_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6535_ net4 mod.des.des_dout\[32\] _3112_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3747_ _0741_ _0742_ _0743_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6466_ _2369_ _3070_ _3074_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3678_ _0663_ _3215_ _0670_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ _2228_ _2332_ _2337_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5512__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _2961_ _3031_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__A3 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ mod.registers.r3\[2\] _2291_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4287__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _2230_ _2244_ _2245_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4079__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4079__B2 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3826__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3826__B2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5846__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4750__I _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4554__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A1 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4609__A3 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3817__B2 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _1381_ _1590_ _1647_ _1387_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xinput10 io_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3601_ _0593_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5742__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4581_ _1299_ _1202_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6690__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6320_ _0740_ _2977_ _2978_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3532_ _0526_ _0527_ _0528_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6251_ _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3463_ _0452_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5491__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ mod.registers.r1\[5\] _2166_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6182_ mod.des.des_dout\[8\] _2876_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3394_ _3236_ _3237_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ _0944_ _2111_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _1911_ _2036_ _2050_ _0001_ _2051_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_69_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3808__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _0997_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _2695_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4917_ _1545_ _1564_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__I _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ mod.registers.r14\[11\] _2654_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _1768_ _1784_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5733__A1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ mod.ldr_hzd\[12\] _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__B1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6518_ _3104_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6449_ _3061_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6533__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4472__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6524__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4550__I2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__B _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ _2525_ _2605_ _2609_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ mod.registers.r11\[4\] _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5486__I _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4702_ _1638_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5682_ mod.registers.r9\[12\] _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4633_ _1235_ _1260_ _1629_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5715__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4564_ _1462_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6303_ _0830_ _2849_ _2967_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3515_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6515__I0 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _1489_ _1221_ _1057_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _2919_ _2921_ _2799_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3446_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4151__B1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6165_ mod.instr\[4\] _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3377_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6586__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _2818_ _1961_ _2090_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__B _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _1911_ _2023_ _2034_ _2035_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5949_ _2694_ _2697_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3909__I _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__S _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5064__C _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4693__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_303 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_314 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_325 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5080__B _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_336 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_347 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_358 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_369 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4445__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A1 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__B1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5173__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3300_ mod.instr_2\[15\] _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__6122__A1 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4280_ _1277_ _0733_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_4_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4684__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6921_ _0081_ net91 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _0012_ net168 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _2585_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _0346_ net147 mod.pc0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3995_ _0966_ _0990_ _0992_ _3222_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ mod.registers.r10\[15\] _2551_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__C _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5665_ _2203_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3962__A3 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1221_ _1223_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5164__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ mod.registers.r8\[0\] _2463_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4547_ _1341_ _1541_ _1542_ _1479_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_2_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__I _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6113__A1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _0857_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6217_ mod.instr\[17\] _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ mod.registers.r9\[0\] _0423_ _0426_ mod.registers.r3\[0\] _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4675__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3722__I0 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6148_ mod.des.des_dout\[0\] _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6079_ mod.pc\[11\] _1747_ _2054_ _2062_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6601__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3374__I _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4115__B1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4666__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4418__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4933__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout142_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__B1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ mod.registers.r1\[5\] _0747_ _0489_ mod.registers.r13\[5\] _0778_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6343__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__B2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1157_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5381_ _2255_ _2308_ _2313_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4332_ _1281_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net210 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6002_ mod.pc\[1\] _2737_ _2710_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _1176_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _0064_ net212 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6624__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3632__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6835_ _0398_ net173 mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3459__I _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6766_ _0332_ net64 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5385__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ mod.registers.r14\[6\] _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6774__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3396__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5717_ _2532_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3396__B2 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _0263_ net101 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _2157_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5137__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5579_ _2431_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4896__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3922__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3369__I _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5128__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4421__C _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A1 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A3 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6647__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__A1 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__I _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4950_ _0713_ _0719_ _1891_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A1 mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4811__B2 mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6797__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3901_ _3139_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4881_ _1862_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3279__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _0186_ net90 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ mod.pc_2\[1\] _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6551_ _0117_ net129 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3763_ mod.registers.r12\[6\] _0503_ _0621_ mod.registers.r15\[6\] _0761_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _2401_ _2391_ _2402_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6482_ _2389_ _3082_ _3084_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3694_ mod.registers.r15\[2\] _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5433_ _2346_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5364_ mod.registers.r3\[8\] _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3550__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3742__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5295_ _2108_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4246_ _1238_ _1239_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3302__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4177_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0381_ net195 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6749_ _0315_ net63 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3917__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4030__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6307__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3541__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3541__B2 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3652__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__I _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4432__B _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3827__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A1 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__B2 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout105_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _1095_ _1096_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _1064_ _1068_ _3187_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4031_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5982_ _2688_ _2076_ _2719_ _2720_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5588__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _1342_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4864_ _0728_ _1860_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _0169_ net82 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3815_ mod.pc_2\[2\] _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _1775_ _1785_ _1788_ _1776_ _1789_ _1777_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_6534_ _3114_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ mod.registers.r4\[7\] _3259_ _3261_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ mod.registers.r15\[6\] _3071_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3677_ _0671_ _0672_ _0673_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6812__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ mod.registers.r4\[11\] _2333_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _1771_ _3028_ _3029_ _3006_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5512__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5347_ _2144_ _2289_ _2293_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5278_ mod.registers.r1\[13\] _2237_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5276__A1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4079__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4229_ _1012_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4517__B _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5200__A1 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5503__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__I _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__A1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5019__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3600_ _0594_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput11 io_in[1] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _1574_ _1575_ _1576_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5742__A2 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3531_ mod.registers.r7\[14\] _0516_ _0518_ mod.registers.r5\[14\] _0529_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6250_ _1831_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3462_ _0456_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6181_ mod.instr\[8\] _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3292__I _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3393_ mod.instr_2\[13\] _3228_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5132_ net12 _2101_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5258__A1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _1078_ _1083_ _1985_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3808__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ _1007_ _1010_ _1011_ _0535_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_84_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__B _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ _2705_ _1983_ _2709_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4233__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5430__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ _1872_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ _2383_ _2653_ _2657_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5981__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _0729_ _1800_ _1814_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ mod.ldr_hzd\[13\] _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__A1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6517_ mod.des.des_dout\[25\] net10 _3088_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3729_ _0725_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3744__B2 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6533__I1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6379_ _2933_ _1828_ _3008_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A1 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3930__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4472__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__I _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5421__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5857__I _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A3 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__I _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6524__I1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__I3 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4463__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout172_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6372__B _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4215__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _2559_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5963__A2 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4604__C _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4701_ _1452_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5681_ _2490_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3287__I _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _1397_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _1052_ _1219_ _1216_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ mod.pc_1\[1\] _2966_ _2964_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3514_ _0425_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6515__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4494_ _1488_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5479__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ _1346_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3445_ _3200_ _3218_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6140__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4151__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ _2865_ _2867_ _2868_ _2859_ _2869_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__B2 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3376_ mod.instr_2\[12\] _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ net11 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6095_ _2784_ _2808_ _2815_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1115_ _1120_ _1985_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _2688_ _1908_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3965__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _2639_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6502__S _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__A3 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3717__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3925__I _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6301__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_304 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_315 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_326 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_337 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_348 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_359 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4445__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3653__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A2 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4705__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6442__I0 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__B2 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6211__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4133__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3570__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5633__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _0080_ net54 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3644__B1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6851_ _0011_ net170 mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _2507_ _2593_ _2598_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6782_ _0345_ net150 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3994_ _0596_ mod.funct3\[1\] _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5733_ _2525_ _2550_ _2554_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _2507_ _2500_ _2508_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4615_ _1228_ _1229_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5595_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4546_ _1462_ _1396_ _1397_ _1031_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6553__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _0737_ _0703_ _1279_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5960__I _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6216_ _2906_ _2903_ _2907_ _2908_ _2905_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3428_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4675__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3722__I1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3359_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6078_ _2784_ _2796_ _2801_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5029_ mod.pc0\[8\] _1905_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3635__B1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6352__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4363__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__I _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4115__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__B2 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5863__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3390__I mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3929__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__B2 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3565__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _1155_ _1260_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5380_ mod.registers.r3\[15\] _2309_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _1313_ _1320_ _1323_ _1325_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout209 net210 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4262_ _0866_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4657__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2724_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5854__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _0914_ _1190_ _0958_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_79_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _0063_ net212 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _0397_ net172 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A1 _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6765_ _0331_ net66 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ _0972_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ _2530_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3396__A2 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _0262_ net106 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _2495_ _2489_ _2496_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _2387_ _2445_ _2450_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4896__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _0736_ _1382_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5690__I _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3305__C1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3608__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6599__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4033__B1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4336__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4639__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 io_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4880_ _1866_ _1875_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3831_ _0600_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6380__B _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6550_ _0116_ net130 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3762_ _0756_ _0757_ _0758_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5501_ mod.registers.r5\[15\] _2392_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ mod.registers.r15\[12\] _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5119__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3693_ mod.registers.r12\[2\] _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _2290_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _0828_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3550__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _2118_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _1241_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3838__B1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3302__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _0544_ _1171_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6817_ _0380_ net195 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4566__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4566__B2 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _0314_ net100 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4030__A3 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _0245_ net101 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4318__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3526__C1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__I _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5818__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__B1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5595__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__S _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6614__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__A2 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4030_ _0535_ _0479_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6764__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _2687_ _2075_ _2078_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _1884_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3599__A2 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4863_ _3195_ _3196_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _0168_ net83 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3814_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4794_ _1774_ _1787_ _0583_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6533_ net3 mod.des.des_dout\[31\] _3112_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3745_ mod.registers.r2\[7\] _0483_ _3254_ mod.registers.r11\[7\] _0743_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _2366_ _3070_ _3073_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3676_ mod.registers.r2\[8\] _0484_ _0415_ mod.registers.r5\[8\] _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5415_ _2221_ _2332_ _2336_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3753__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _2961_ _3030_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3523__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ mod.registers.r3\[1\] _2291_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6473__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _0997_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _0561_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3928__I _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6637__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4711__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__B2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 io_in[2] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout215_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3530_ mod.registers.r2\[14\] _0485_ _0513_ mod.registers.r3\[14\] _0528_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4950__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3461_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ mod.des.des_dout\[26\] _2151_ _2170_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6180_ _2878_ _2879_ _2880_ _2872_ _2881_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3392_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ mod.valid2 _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _2037_ _2039_ _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4013_ _0448_ mod.funct3\[0\] _0886_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__B2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2706_ mod.pc0\[6\] _2707_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5430__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _1873_ _1894_ _1909_ _1910_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3441__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ mod.registers.r14\[10\] _2654_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5981__A3 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3992__A2 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4846_ _0729_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ mod.ldr_hzd\[14\] _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6516_ _3103_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ _0446_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6447_ _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3659_ mod.registers.r9\[9\] _0623_ _0624_ mod.registers.r3\[9\] _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5497__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1767_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _2262_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6446__A1 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A4 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3983__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout165_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3568__I _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4700_ _0767_ _1018_ _1611_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5680_ _2488_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4631_ _1235_ _1434_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3726__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _1281_ _1551_ _1553_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6301_ _2678_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3513_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4493_ _1014_ _1490_ _1015_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6232_ _2678_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3444_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ _2683_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3375_ mod.instr_2\[13\] _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _2095_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout78_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ mod.pc\[13\] _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ _1895_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__B _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5947_ _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3478__I _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _2358_ _2640_ _2646_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5167__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ _1816_ _1817_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4509__A4 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_305 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4258__B _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_316 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_327 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_338 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6029__I mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_349 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3653__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5868__I _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3653__B2 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__I mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6442__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A2 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3337__B _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5330__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__B1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5633__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3644__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3644__B2 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__B1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6850_ _0010_ net168 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ mod.registers.r12\[7\] _2594_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5397__A1 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _0344_ net150 mod.pc0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4444__I0 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3993_ _0886_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5732_ mod.registers.r10\[14\] _2551_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5663_ mod.registers.r9\[7\] _2501_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__I _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _1610_ _1016_ _1488_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5594_ _2459_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4545_ _1029_ _1500_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5018__I _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4476_ _1451_ _1472_ _1341_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6215_ _1856_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5321__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ _3249_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6848__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3332__B1 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__A3 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6146_ _2673_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ _3209_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _2737_ _2802_ _2803_ _2719_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3289_ _3136_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _2008_ _2016_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3635__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3635__B2 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6424__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6513__S _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3936__I _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4363__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5312__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5863__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6040__A2 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout128_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ _1326_ _1327_ _1273_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5303__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0861_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _2729_ _2735_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5854__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _1185_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input2_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__B _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ _0062_ net215 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4345__C _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6833_ _0396_ net172 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _0330_ net100 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3976_ _3173_ _0580_ mod.registers.r1\[6\] _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5715_ _2507_ _2538_ _2543_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5790__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _0261_ net101 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ mod.registers.r9\[2\] _2491_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5542__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5577_ mod.registers.r7\[11\] _2446_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _1438_ _0677_ _1379_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4459_ _1454_ _1455_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3491__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3305__B1 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5845__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3305__C2 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3856__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ mod.pc_1\[9\] _2841_ _2837_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3608__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3608__B2 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5211__I _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4033__B2 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6418__S _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__I mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ _0738_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5221__B1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__A1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ mod.registers.r4\[6\] _0638_ _3262_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3576__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6693__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6480_ _3064_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3692_ _3175_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5431_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5524__A1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3535__B1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5362_ _2288_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _1283_ _1294_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _2113_ _2116_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0662_ _1121_ _1123_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3838__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3838__B2 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4175_ _1172_ _1156_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5966__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _0379_ net153 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4015__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4566__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _0313_ net63 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3959_ _0953_ _0954_ _0955_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3486__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3774__B1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _0244_ net105 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _2395_ _2480_ _2483_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5515__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__B1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__C2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4629__I0 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__B2 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4557__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5754__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__B1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4309__A2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4020__I _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5809__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6909__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__A2 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout195_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4176__B _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3679__S0 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _1911_ _1913_ _1924_ _1925_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6391__B _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _1857_ _1858_ _1859_ _1348_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _0167_ net126 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ _0799_ _3262_ _0804_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5745__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _1786_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6532_ _3113_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3744_ mod.registers.r6\[7\] _0634_ _0491_ mod.registers.r14\[7\] _0742_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6463_ mod.registers.r15\[5\] _3071_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3675_ mod.registers.r9\[8\] _0623_ _0605_ mod.registers.r14\[8\] _0673_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5414_ mod.registers.r4\[10\] _2333_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _1772_ _3028_ _3029_ _1828_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3603__S0 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5345_ _2135_ _2289_ _2292_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3523__A3 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4720__A2 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6589__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5276_ mod.des.des_dout\[34\] _2171_ _2240_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ _0994_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6473__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4158_ _1154_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4086__B _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4089_ _0463_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5736__A1 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3598__I0 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__B1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6464__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4724__B _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6431__S _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[3] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3854__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4950__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout110_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout208_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3460_ _0457_ _0450_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _3241_ _3242_ _3236_ _3237_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _2109_ _1848_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _1980_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6881__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ _3221_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _2705_ _1963_ _2708_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ _3188_ _1049_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5894_ _2380_ _2653_ _2656_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5718__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _1835_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3992__A3 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4776_ mod.ldr_hzd\[15\] _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6515_ mod.des.des_dout\[24\] net9 _3099_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3727_ _3199_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _2286_ _2583_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3658_ mod.registers.r7\[9\] _0418_ _0415_ mod.registers.r5\[9\] _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ _3002_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ _0585_ _0586_ mod.registers.r14\[1\] _0582_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5328_ _2260_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__B _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6315__I _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6604__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3432__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3983__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4448__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout190 net191 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout158_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A3 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ _1627_ _1597_ _1438_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5176__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _1380_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3726__A3 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6300_ _3224_ _2849_ _2965_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3512_ _0430_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4492_ _1034_ _1053_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6231_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3443_ _3199_ _3201_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4687__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4687__B2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6162_ mod.des.des_dout\[3\] _2863_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _3225_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3533__B _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5113_ _1347_ net22 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6093_ _2725_ _2816_ _2817_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _1882_ _2030_ _2031_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6627__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _2096_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ mod.registers.r14\[3\] _2642_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5167__A2 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5195__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4914__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ net13 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6116__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ mod.des.des_dout\[5\] net3 _3050_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3350__A1 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_306 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_317 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_328 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_339 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6107__A1 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__B1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3644__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__B2 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3579__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ _2505_ _2593_ _2597_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _0343_ net150 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5397__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3992_ _0442_ _0970_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4444__I1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ _2523_ _2550_ _2553_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5794__I _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6346__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _2194_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _1016_ _1488_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4544_ _1289_ _1293_ _1313_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1204_ _1451_ _1472_ _1418_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ mod.des.des_dout\[16\] _2900_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout90_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3426_ _3252_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5321__A2 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3332__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ mod.instr\[0\] _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3332__B2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3357_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ mod.pc\[10\] _2724_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3288_ mod.registers.r7\[0\] _3135_ _3139_ mod.registers.r3\[0\] _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6066__S _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _1989_ _2006_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3635__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3489__I _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _1746_ _1849_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4060__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6337__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4113__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3323__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3874__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5879__I _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3399__I _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _0875_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4191_ _1186_ _1187_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _0061_ net215 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0395_ net172 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _0329_ net58 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ _3141_ _3180_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5714_ mod.registers.r10\[7\] _2539_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _0260_ net105 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5790__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _2148_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _2384_ _2445_ _2449_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5542__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3553__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _1312_ _0798_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4868__I _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4458_ _0781_ _1227_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3305__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3409_ _3219_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3305__B2 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4389_ _1279_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _2787_ _2840_ _2842_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ _2787_ _2018_ _1960_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3608__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6524__S _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4033__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3792__B2 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__I _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3847__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__B _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5221__A1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ mod.registers.r2\[6\] _0484_ _3255_ mod.registers.r11\[6\] _0758_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _3171_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _2120_ _2315_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5524__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3535__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _2195_ _2296_ _2301_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _1296_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5292_ _2230_ _2255_ _2256_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5288__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _1240_ _1124_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3838__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4174_ _1142_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3471__B1 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _0378_ net152 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4015__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__C _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6746_ _0312_ net67 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5763__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ mod.registers.r7\[7\] _0679_ _0690_ mod.registers.r14\[7\] _0956_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3774__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6677_ _0243_ net131 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3889_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ mod.registers.r8\[13\] _2481_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5515__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__A1 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__B2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ _2431_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6318__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4629__I1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4254__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A3 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__B2 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4565__I0 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6002__B _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4301__I _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4190__B2 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6429__S _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3296__A3 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout188_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3679__S1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _1891_ _1030_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _0874_ _1739_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6600_ _0166_ net127 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3812_ _0805_ _0806_ _0807_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5745__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _1764_ _1787_ _1788_ _1766_ _1789_ _1767_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3756__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ mod.registers.r8\[7\] _3233_ _0632_ mod.registers.r10\[7\] _0741_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6531_ net2 mod.des.des_dout\[30\] _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3674_ mod.registers.r10\[8\] _0602_ _0627_ mod.registers.r13\[8\] _0672_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6462_ _2361_ _3070_ _3072_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4556__I0 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5413_ _2214_ _2332_ _2335_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6393_ _2104_ _2932_ _2992_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3603__S1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4211__I mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ mod.registers.r3\[0\] _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4181__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _2155_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4226_ _0964_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4484__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__I _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _1142_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _0616_ _0991_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__I _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__C _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__B2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3497__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3598__I1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _0295_ net115 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3762__A4 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5672__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__B1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4791__I _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 io_in[4] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout103_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__B2 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3390_ mod.instr_2\[12\] _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _2040_ _2036_ _2045_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4466__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ _0696_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5663__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3674__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _2706_ mod.pc0\[5\] _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _1895_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5893_ mod.registers.r14\[9\] _2654_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3441__A3 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4206__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ mod.instr_2\[6\] _1838_ _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3729__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _1769_ _1770_ _1771_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6514_ _3102_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3726_ _0500_ _0505_ _0509_ _0520_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6445_ _3060_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3657_ _0651_ _0652_ _0653_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6143__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3588_ _3147_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6376_ _3014_ _3016_ _3010_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__I _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5327_ _2228_ _2274_ _2279_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5258_ mod.des.des_dout\[32\] _2207_ _2224_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ _0732_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5189_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5406__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__I _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3432__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6134__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4145__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout180 net181 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net197 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4081__B1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6442__S _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A4 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4384__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ _1265_ _1556_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3511_ mod.registers.r9\[15\] _0507_ _0508_ mod.registers.r10\[15\] _0509_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4491_ _1058_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3442_ _3224_ _3226_ _0410_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6230_ _2668_ _2681_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5884__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3373_ _3220_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _2094_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6092_ mod.pc\[12\] _2730_ _2812_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4439__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5043_ mod.pc\[9\] _1875_ _1748_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__B1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6061__A1 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5945_ _2685_ mod.pc0\[2\] _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _2355_ _2640_ _2645_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4827_ _1821_ _1817_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4758_ _1752_ _1344_ _1753_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ mod.registers.r7\[4\] _0679_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__I mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _0737_ _1620_ _1686_ _1203_ _1279_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_107_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4127__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6428_ _3051_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4678__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5875__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ _3002_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3350__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_307 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_318 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_329 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4835__C1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4063__B1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4290__B _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4118__B2 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4669__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5094__A2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout170_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _0975_ _0981_ _0985_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4444__I2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ mod.registers.r10\[13\] _2551_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5661_ _2505_ _2500_ _2506_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6346__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _1225_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5592_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _1462_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4109__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4474_ _1459_ _1471_ _1409_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ mod.instr\[16\] _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3425_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__A2 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _3192_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6144_ _2818_ _2851_ _2853_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6075_ _2797_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3287_ _3138_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6282__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _2012_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6146__I _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__A1 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__B1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4596__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ mod.valid1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6894__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _2389_ _2632_ _2634_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6337__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5848__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6025__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4587__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6617__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3364__B _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4511__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ mod.registers.r6\[14\] _0903_ _0920_ mod.registers.r15\[14\] _1188_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6767__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _0060_ net214 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6831_ _0394_ net173 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__D _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _0328_ net67 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3974_ _0476_ _0971_ mod.registers.r8\[6\] _0581_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5713_ _2505_ _2538_ _2542_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6693_ _0259_ net131 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5644_ _2493_ _2489_ _2494_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5575_ mod.registers.r7\[10\] _2446_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ _1489_ _1396_ _1260_ _1057_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _1390_ _1383_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4502__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3305__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3408_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4388_ _1382_ _1384_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3856__A3 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ mod.pc_1\[8\] _2841_ _2837_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ mod.funct3\[2\] _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__A1 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6058_ mod.pc\[8\] _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5009_ _1947_ _1948_ _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__B2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3449__B _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3792__A2 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6246__A1 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout133_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ mod.registers.r11\[2\] _0577_ _0574_ mod.registers.r8\[2\] _0688_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3535__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ mod.registers.r3\[7\] _2297_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4311_ _1285_ _1303_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ mod.registers.r1\[15\] _2237_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4242_ _1111_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3299__A1 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4591__S0 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4637__C _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__I _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A1 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3471__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__B2 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6814_ _0377_ net153 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6745_ _0311_ net102 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3957_ mod.registers.r3\[7\] _0680_ _3144_ mod.registers.r4\[7\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4971__A1 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3774__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _0242_ net121 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3888_ _0726_ _0441_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6932__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ _2390_ _2480_ _2482_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3783__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3526__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _2359_ _2432_ _2438_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _0884_ _0723_ _1379_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5489_ mod.registers.r5\[12\] _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5279__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6535__S _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3462__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__B2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3765__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4789__I _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__I mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4190__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__B _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6219__B2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A3 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _1351_ _1736_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3811_ mod.registers.r1\[3\] _0430_ _0432_ mod.registers.r13\[3\] _0808_ _0809_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ _3178_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _3105_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3756__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3742_ mod.pc_2\[7\] _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4953__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ mod.registers.r15\[4\] _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3673_ mod.registers.r1\[8\] _0510_ _0624_ mod.registers.r3\[8\] _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4705__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ mod.registers.r4\[9\] _2333_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4556__I1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6392_ _3002_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5343_ _2290_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6458__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _2009_ _2129_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _1014_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5130__A1 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _0586_ _1050_ _0934_ _0935_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_110_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _0991_ _1008_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5993__I _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _0294_ net117 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6659_ _0225_ net115 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5672__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3683__B2 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5424__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3688__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput15 io_in[5] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A2 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__B _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5143__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _0889_ mod.funct7\[1\] _0595_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3674__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__B2 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__C _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _2695_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4912_ _1749_ _1904_ _1906_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ _2375_ _2653_ _2655_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5179__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4843_ _1839_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4931__B _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3729__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ mod.ldr_hzd\[8\] _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6513_ mod.des.des_dout\[23\] net8 _3099_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3725_ _0705_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5318__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ mod.des.des_dout\[12\] net10 _3044_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3656_ mod.registers.r4\[9\] _3260_ _3221_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A1 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _2999_ _3015_ _3008_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3587_ _3181_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5326_ mod.registers.r2\[11\] _2275_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6149__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _2124_ _2225_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ _1200_ _1201_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5188_ mod.des.des_dout\[25\] _2125_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4139_ _1074_ _1134_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5893__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3656__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout181 net182 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout192 net196 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4081__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4081__B2 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5581__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout213_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3510_ _3239_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4490_ _1487_ _1455_ _1453_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4977__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A1 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3441_ _0416_ _0419_ _0427_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_109_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5884__A2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _2673_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ mod.pc_2\[0\] _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5111_ _1760_ _1849_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _2809_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ mod.pc0\[9\] _1905_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3647__B2 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6436__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5944_ _2693_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4072__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ mod.registers.r14\[2\] _2642_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4826_ _1781_ _1820_ _1823_ _1779_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1752_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6673__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _0441_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4688_ _0884_ _1506_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6427_ mod.des.des_dout\[4\] net2 _3050_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3639_ mod.registers.r2\[10\] _3251_ _0636_ mod.registers.r11\[10\] _0637_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6358_ _2698_ _1763_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__C _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5309_ _2262_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _2955_ _2958_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_308 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_319 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__B1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__C2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6543__S _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4063__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4063__B2 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3810__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3810__B2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4366__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5315__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4746__B _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__B1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6418__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6546__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout163_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _0986_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4444__I3 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__I _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ mod.registers.r9\[6\] _2501_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4611_ _3217_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5554__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5591_ _2316_ _2458_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _1539_ _1023_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5306__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4109__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _1464_ _1469_ _1470_ _1222_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6212_ _2902_ _2903_ _2904_ _2896_ _2905_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3317__B1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3424_ _0420_ _0421_ _0412_ _0413_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__3868__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ mod.pc_1\[13\] _2852_ _2844_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3355_ _3206_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2049_ _2800_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__B _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3286_ _3133_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5025_ _2013_ _1996_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__B2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ mod.registers.r13\[12\] _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5545__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _1802_ _0429_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5789_ mod.registers.r12\[2\] _2588_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3556__B1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5506__I _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4410__I _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5839__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3364__C _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__B _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6247__I _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0393_ net173 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5775__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4578__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _0327_ net100 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3973_ _3130_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5712_ mod.registers.r10\[6\] _2539_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _0258_ net120 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5643_ mod.registers.r9\[1\] _2491_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _2381_ _2445_ _2448_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4525_ _1055_ _0861_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6711__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4387_ _1265_ _0601_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _2826_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3710__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _3124_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _2779_ _2786_ _2684_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3269_ mod.des.des_counter\[0\] _3120_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6861__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5008_ _1989_ _1997_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4018__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3777__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__C mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3529__B1 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5236__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4140__I mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4009__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3480__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4315__I _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3768__B1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5509__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6530__I _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6734__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4050__I _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4310_ _1304_ _1305_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4241_ _1108_ _1109_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _0982_ _1050_ _0934_ _0935_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_67_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4591__S1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4248__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5996__A1 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A2 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _0376_ net159 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout39_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3759__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3956_ mod.registers.r1\[7\] _3149_ _3168_ mod.registers.r8\[7\] _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6744_ _0310_ net104 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _0241_ net132 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4971__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3887_ _3159_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5626_ mod.registers.r8\[12\] _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4184__B1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__A1 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ mod.registers.r7\[3\] _2434_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4508_ _1266_ _0702_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _2349_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6476__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _1207_ _1277_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6228__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _2811_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6607__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__B2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4714__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5978__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _0471_ _3231_ _0435_ _0436_ _0472_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4790_ _0982_ _0445_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3741_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _3064_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3672_ _0664_ _0665_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4166__B1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5411_ _2204_ _2332_ _2334_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5902__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6391_ _3025_ _3027_ _3022_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__B1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5342_ _2287_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6458__A2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _1209_ _2152_ _2172_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4469__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__C _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4224_ _1055_ _1056_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _1048_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5969__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4086_ _0706_ _1078_ _1083_ _0966_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_37_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6435__I _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6394__A1 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__B2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _1960_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6727_ _0293_ net104 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3939_ _0881_ _0891_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4944__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3747__A3 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _0224_ net112 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _2367_ _2468_ _2471_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6589_ _0155_ net81 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A3 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3994__I0 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 io_in[6] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__B1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4699__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout193_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _2698_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4911_ mod.pc\[2\] _1865_ _1867_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5891_ mod.registers.r14\[8\] _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5179__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4842_ _1770_ _1825_ _1827_ _1772_ mod.instr_2\[5\] _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4931__C _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ mod.ldr_hzd\[9\] _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4503__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _3101_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3724_ _0706_ _0713_ _0719_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__6128__A1 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _3059_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3655_ mod.registers.r2\[9\] _0484_ _3255_ mod.registers.r11\[9\] _0653_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6374_ _1823_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3586_ mod.registers.r12\[1\] _0581_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5325_ _2221_ _2274_ _2278_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__C _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5256_ _1969_ _2181_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6300__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5187_ _2161_ _2127_ _2132_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4862__B2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _1135_ _1069_ _1071_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__I mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input19_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4069_ mod.registers.r6\[11\] _0902_ _0928_ mod.registers.r13\[11\] _1067_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__B1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A2 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6119__A1 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout160 net161 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout171 net174 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3656__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout182 net198 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout193 net196 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3699__I _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5419__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A1 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3592__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3440_ mod.registers.r1\[0\] _0431_ _0433_ mod.registers.r13\[0\] _0437_ _0438_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_fanout206_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3371_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _1945_ _1190_ _2093_ _1873_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ _2814_ _2077_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _2008_ _2028_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4993__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3647__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3402__I _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _0003_ _2691_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _2352_ _2640_ _2644_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__I _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5572__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ mod.pc_2\[0\] _1011_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ _3226_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _1325_ _1368_ _1652_ _1439_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6426_ _3044_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3638_ _3254_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5324__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6357_ _2104_ _2671_ _3001_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3569_ mod.registers.r4\[1\] _0565_ _0566_ mod.registers.r1\[1\] _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5308_ _2260_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _0476_ _2957_ _2953_ mod.instr\[17\] _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_309 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _2154_ _2023_ _2208_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4835__A1 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__B2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4063__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5012__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5563__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__B1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5079__A1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4054__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout156_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__B1 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _1538_ _1545_ _1564_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5590_ _2103_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4541_ _1465_ _1467_ _1468_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4988__I _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ _1224_ _1225_ _1014_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3317__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6211_ _2718_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3423_ _3228_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3317__B2 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _2826_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3354_ _3193_ _3198_ _3205_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _1346_ _1746_ _2038_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3285_ _3136_ mod.instr_2\[16\] _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1990_ _1993_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5490__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4228__I _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__A1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6640__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _2614_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4808_ mod.ldr_hzd\[8\] _0434_ _0616_ _0615_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5545__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _2493_ _2586_ _2590_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3556__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3556__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _1351_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4505__B1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _3038_ _3039_ _2732_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__I _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3795__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3547__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5432__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5472__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6663__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ _0326_ net103 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _0967_ _0968_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ _2503_ _2538_ _2541_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3786__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _0257_ net120 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ _2143_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3538__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3836__B _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ mod.registers.r7\[9\] _2446_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _1418_ _1496_ _1504_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _0780_ _1012_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3406_ _3241_ _3257_ _3231_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4386_ _1383_ _1354_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3710__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _3151_ _3186_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6125_ _2670_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3710__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _2000_ _2780_ _2781_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_85_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3268_ _3122_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _1896_ _1988_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3797__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3777__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5909_ net11 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6889_ _0049_ net166 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3746__B _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__B2 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5517__I _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4257__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4009__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3500__I _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3768__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3768__B2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5509__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3656__B _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4568__I0 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4193__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1128_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4171_ _1048_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4248__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _0375_ net159 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3410__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A2 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3759__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3759__B2 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6743_ _0309_ net103 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__B _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3955_ mod.registers.r12\[7\] _0716_ _0689_ mod.registers.r13\[7\] _0953_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6674_ _0240_ net132 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3886_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ _2462_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4184__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _2356_ _2432_ _2437_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4507_ _0938_ _1383_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5487_ _2347_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _1366_ _1435_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _1172_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3695__B1 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _1879_ _2825_ _2829_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4239__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _2761_ _2763_ _1956_ _2769_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3998__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6539__I1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4175__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5427__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3989__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _0464_ _0700_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4953__A3 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _3202_ _0666_ _0667_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ mod.registers.r4\[8\] _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6851__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4166__B2 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _3026_ _3015_ _3007_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5902__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3913__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5341_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3913__B2 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5272_ _2140_ _2081_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5106__B _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ _1216_ _1217_ _1219_ _1220_ _1029_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4154_ _1147_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4085_ _1079_ _1080_ _1081_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3429__B1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout51_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4236__I _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ mod.pc0\[6\] _1958_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6726_ _0292_ net106 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3938_ _0913_ _0933_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3747__A4 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6657_ _0223_ net38 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3869_ _0457_ _0456_ _0451_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4157__A1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ mod.registers.r8\[5\] _2469_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6588_ _0154_ net81 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5539_ _2390_ _2424_ _2426_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5657__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__B1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__I1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 io_in[7] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4148__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__B2 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__B1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A2 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout186_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__C _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__B1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ mod.pc0\[2\] _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5890_ _2641_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4841_ _1771_ _1820_ _1823_ _1769_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3895__I _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5088__S _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4387__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4772_ mod.ldr_hzd\[10\] _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6511_ mod.des.des_dout\[22\] net7 _3099_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3723_ _0444_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6128__A2 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6442_ mod.des.des_dout\[11\] net9 _3055_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3654_ mod.registers.r8\[9\] _3234_ _0602_ mod.registers.r10\[9\] _0652_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5887__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _1779_ _3003_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5615__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3585_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4659__C _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ mod.registers.r2\[10\] _2275_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout99_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5255_ _2127_ _2053_ _2208_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6300__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5186_ _2126_ _1928_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _0631_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ mod.registers.r11\[11\] _0916_ _0925_ mod.registers.r1\[11\] _1066_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4614__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5811__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6897__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__B1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__I mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__B2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _0275_ net133 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout150 net154 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout161 net162 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout172 net174 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout183 net186 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout194 net196 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5802__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__B1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6305__B _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3592__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout101_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ _3221_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _1989_ _2023_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__B _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5942_ _2690_ mod.pc0\[1\] _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3804__B1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ mod.registers.r14\[1\] _2642_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _1821_ _1818_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5021__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ mod.pc_2\[0\] _1011_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3706_ _0482_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4780__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _1180_ _1370_ _1546_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6425_ _3049_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3637_ mod.registers.r6\[10\] _0634_ _3247_ mod.registers.r14\[10\] _0635_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4532__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ mod.rd_3\[3\] _2824_ _2097_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3568_ _3148_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _2158_ _2261_ _2267_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ _2934_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3499_ _3255_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5238_ _2024_ _2198_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__I mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _2139_ _1894_ _2132_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4048__B1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3271__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3810__A3 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__B _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6912__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__B2 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5079__A2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6086__I _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3503__I _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout149_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__B2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _1524_ _1531_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4762__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6592__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _1465_ _1467_ _1468_ _1461_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5165__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ mod.des.des_dout\[15\] _2900_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3422_ _3227_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3317__A2 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2670_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _3204_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2791_ _2798_ _2799_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3284_ mod.instr_2\[17\] _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _1990_ _1993_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5242__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _2676_ _1847_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5856_ _2612_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6935__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ _1782_ mod.ldr_hzd\[1\] mod.ldr_hzd\[2\] mod.ldr_hzd\[3\] _1801_ _1802_ _1805_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5787_ mod.registers.r12\[1\] _2588_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3556__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4753__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _1715_ _1735_ _1518_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3800__I0 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _1420_ _1661_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6408_ _3026_ _3006_ _3036_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6339_ _2111_ _2990_ _2799_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5803__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A1 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3795__A2 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3547__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3952__C1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6249__A1 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3971_ mod.registers.r11\[6\] _3166_ _0578_ mod.registers.r10\[6\] mod.registers.r2\[6\]
+ _0922_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_16_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ mod.registers.r10\[5\] _2539_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3786__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _0256_ net131 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5641_ _2486_ _2489_ _2492_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4999__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5572_ _2376_ _2445_ _2447_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _3209_ _1492_ _1517_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3408__I _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4454_ _1224_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ _3242_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _1276_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6124_ _2001_ _2833_ _2839_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3710__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _1882_ _1876_ _2784_ _2687_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3267_ net184 _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _1990_ _1993_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_54_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _2400_ _2659_ _2664_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3777__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6888_ _0048_ net166 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5839_ _2361_ _2620_ _2622_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3529__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__S0 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3701__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4257__A3 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5206__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3768__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3937__B _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4612__I _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4568__I1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5390__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4193__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__C _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _1160_ _1161_ _1162_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6493__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6780__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3456__A1 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3898__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ _0374_ net159 mod.pc_1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6742_ _0308_ net103 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3759__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ _0949_ _0950_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6673_ _0239_ net38 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3885_ _0881_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4522__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5624_ _2460_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4184__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5381__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ mod.registers.r7\[2\] _2434_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _1454_ _1258_ _1499_ _1375_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5133__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _0882_ _0797_ _0702_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5353__I _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4368_ _1271_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ mod.pc_1\[1\] _2827_ _2812_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3319_ _3145_ _3147_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ mod.pc_2\[7\] _1176_ _0745_ _0753_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ _2768_ _2764_ _1956_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6359__I _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5675__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__B _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6094__I mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3989__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6027__C _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__I _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout131_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3670_ _0612_ _0616_ mod.registers.r8\[8\] _0610_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5271_ _2230_ _2236_ _2238_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ _1047_ _1051_ _1029_ _1031_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_68_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ _1148_ _1149_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ mod.registers.r5\[10\] _0568_ _0565_ mod.registers.r4\[10\] _1082_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3429__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3429__B2 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_290 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout44_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _1853_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6725_ _0291_ net134 mod.registers.r12\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _0889_ _0934_ _0725_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3601__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _0222_ net39 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ _0865_ _3206_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _2362_ _2468_ _2470_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4157__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5354__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _0153_ net81 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3799_ _0599_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5538_ mod.registers.r6\[12\] _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _2347_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3380__A3 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5967__B _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3840__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__B2 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 io_in[8] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5345__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A2 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__I _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__B2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6549__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__B _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout179_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4084__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3831__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6699__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _1831_ _1836_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4387__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ mod.ldr_hzd\[11\] _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _3100_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3722_ mod.funct7\[1\] mod.funct7\[0\] _0595_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4792__C1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _3058_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5336__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3653_ mod.registers.r6\[9\] _0604_ _0605_ mod.registers.r14\[9\] _0651_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5887__A2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ _3011_ _3013_ _3010_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3584_ _3136_ _3162_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5323_ _2214_ _2274_ _2277_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5254_ _2057_ _2198_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ mod.pc_2\[4\] _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4136_ _1128_ _1131_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ mod.registers.r14\[11\] _0917_ _0930_ mod.registers.r9\[11\] mod.registers.r2\[11\]
+ _0923_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4075__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__A1 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__B2 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _1957_ _1854_ _1959_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6708_ _0274_ net120 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5327__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _0205_ net51 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5878__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3326__I _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout151 net153 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout162 net199 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout173 net174 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout184 net186 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout195 net196 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6841__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5716__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6046__A2 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _1881_ _1889_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3804__B2 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _2344_ _2640_ _2643_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4823_ _1816_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5557__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__S _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4754_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3705_ _0601_ _0677_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _1211_ _1370_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4780__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ mod.des.des_dout\[3\] net19 _3045_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3636_ _3243_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _2999_ _2671_ _3000_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4532__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3567_ _3143_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5306_ mod.registers.r2\[3\] _2263_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6286_ _2955_ _2956_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4686__B _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3498_ mod.registers.r13\[15\] _0490_ _0492_ mod.registers.r14\[15\] mod.registers.r15\[15\]
+ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6285__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ _2181_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6864__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _1897_ _2140_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ mod.registers.r5\[9\] _0897_ _0899_ mod.registers.r3\[9\] _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5099_ mod.pc\[13\] _1876_ _1867_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A1 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4048__B2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__B _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__I mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3271__A2 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3559__B1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__I _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__I _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__I _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6737__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5446__I _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout211_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__I _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3970__B1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1047_ _1051_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ mod.registers.r7\[0\] _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2847_ _2849_ _2850_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _2666_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5181__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4278__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _2010_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3789__B1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5924_ net12 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5855_ _2386_ _2626_ _2631_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _0615_ _0607_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4202__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _2486_ _2586_ _2589_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4737_ _1337_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4753__A2 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4260__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3800__I1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4668_ _1663_ _1665_ _1609_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4505__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3619_ _0428_ _0609_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6407_ _1776_ _3034_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _1596_ _0460_ _0846_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ mod.valid_out3 _2112_ _2848_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _2941_ _2945_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5975__B _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__A1 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3952__C2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3514__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3450__S _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__I0 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout161_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ mod.registers.r5\[6\] _0896_ _0575_ mod.registers.r9\[6\] _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4432__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ mod.registers.r9\[0\] _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5571_ mod.registers.r7\[8\] _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4522_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A2 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4453_ _1022_ _1059_ _1239_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3404_ mod.registers.r2\[0\] _3251_ _3255_ mod.registers.r11\[0\] _3256_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4384_ _0882_ _0702_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ mod.pc_1\[7\] _2834_ _2837_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3335_ _3123_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5999__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3266_ _0000_ _3120_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4120__B1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5005_ _1994_ _1972_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ mod.registers.r14\[15\] _2660_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6887_ _0047_ net167 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6470__I _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ mod.registers.r13\[4\] _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _2557_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3934__B1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__I _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6582__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4009__A4 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3509__I _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5390__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__B1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3456__A2 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__I0 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6491__S _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6810_ _0373_ net187 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _0307_ net116 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4956__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3953_ mod.registers.r2\[7\] _0922_ _3166_ mod.registers.r11\[7\] _0951_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6158__B2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3884_ _0521_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6672_ _0238_ net38 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4169__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5905__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _2387_ _2474_ _2479_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5554_ _2353_ _2432_ _2436_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4505_ _1228_ _1259_ _1501_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5485_ _2235_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5634__I _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5133__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _1361_ _1364_ _1304_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3695__A2 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _2727_ _2825_ _2828_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3318_ _3136_ _3162_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4298_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6037_ _1345_ _1745_ _1957_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4644__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _0099_ net213 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4947__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4635__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__C _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A3 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6388__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__C _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ mod.registers.r1\[12\] _2237_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4221_ _1218_ _0867_ _1037_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4152_ mod.registers.r5\[12\] _0898_ _0920_ mod.registers.r15\[12\] _1150_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4083_ mod.registers.r7\[10\] _0679_ _0710_ mod.registers.r15\[10\] _1081_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3429__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_280 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4019__B _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_291 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6379__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ mod.pc\[6\] _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5051__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _0290_ net121 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3936_ _3218_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3601__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ _0221_ net53 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ _0850_ _0852_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5606_ mod.registers.r8\[4\] _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6586_ _0152_ net80 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3798_ _0562_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5537_ _2406_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _2375_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4419_ _1355_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5399_ _2320_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3668__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__B _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6620__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 io_in[9] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3659__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__I _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5584__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _1764_ _1765_ _1766_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _0714_ _0717_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4792__B1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__C2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ mod.des.des_dout\[10\] net8 _3055_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3652_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5184__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6371_ _2999_ _3012_ _3008_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3583_ _3181_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5322_ mod.registers.r2\[9\] _2275_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _2197_ _2221_ _2222_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5912__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4847__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _0728_ _0731_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ _2122_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _1132_ _1084_ _1087_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ _1060_ _1061_ _1062_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4075__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6643__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__I _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5575__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3586__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ _0273_ net120 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6793__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _3176_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4899_ _3125_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6638_ _0204_ net51 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5327__A2 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3607__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _0135_ net129 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout130 net136 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout152 net153 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout163 net199 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout174 net181 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3342__I mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout185 net186 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout196 net197 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__A2 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5269__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5015__A1 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4173__I _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4901__I mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4526__B1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5218__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4549__S _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3501__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3501__B2 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout191_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5254__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5940_ _2676_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__A2 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ mod.registers.r14\[0\] _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4753_ _1750_ _1742_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3704_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4684_ _1680_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4780__A3 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6423_ _3048_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3635_ mod.registers.r8\[10\] _0486_ _0632_ mod.registers.r10\[10\] _0633_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6354_ mod.rd_3\[2\] _2824_ _2097_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _0441_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5305_ _2149_ _2261_ _2266_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3740__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6285_ _0697_ _2950_ _2953_ mod.instr\[16\] _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3497_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _2105_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _2123_ _2144_ _2145_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ mod.registers.r10\[9\] _0894_ _0930_ mod.registers.r9\[9\] _1116_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ mod.pc0\[13\] _1978_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4048__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _3226_ _0700_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3559__B2 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4220__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3731__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6689__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A3 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__I _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5787__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4598__I0 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5727__I _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3970__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__B2 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout204_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5711__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _2792_ _2795_ _2797_ _2730_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3282_ _3128_ _3130_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6511__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5475__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _0663_ _2009_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__A3 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__C _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5923_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5854_ mod.registers.r13\[11\] _2627_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _1777_ _1776_ mod.ldr_hzd\[14\] _1774_ _1801_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5785_ mod.registers.r12\[0\] _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5637__I _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _1719_ _1722_ _1723_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3800__I2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3961__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _1252_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _3035_ _3037_ _3022_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3618_ _3257_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0842_ _0825_ _0563_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6337_ _1209_ _2920_ _2989_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5372__I _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3549_ _0545_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ _1801_ _2943_ _2938_ mod.instr\[10\] _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6502__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5466__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _1898_ _2172_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6199_ _1856_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A2 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3952__B2 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__B _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5457__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__B1 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5209__A1 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__B _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout154_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6854__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2433_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3943__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4521_ _0945_ _1518_ _0854_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _1449_ _1414_ _1207_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3403_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _1977_ _2833_ _2838_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _3157_ _3164_ _3169_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2739_ _2755_ _2771_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ mod.des.des_counter\[1\] _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _1968_ _1969_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4120__B2 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout67_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _2397_ _2659_ _2663_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _0046_ net166 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ _2614_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ _2517_ _2571_ _2576_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3934__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3934__B2 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1133_ _1716_ _1245_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _2486_ _2531_ _2534_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5439__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__B _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4717__A3 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3689__B1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5740__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__B2 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__B _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3456__A3 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4356__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3700__I1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _0306_ net115 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3952_ mod.registers.r15\[7\] _0589_ _0711_ mod.registers.r9\[7\] mod.registers.r6\[7\]
+ _0572_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _0237_ net53 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6158__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4305__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3883_ _0853_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4169__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ mod.registers.r8\[11\] _2475_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5905__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ mod.registers.r7\[1\] _2434_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1226_ _1227_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5484_ _2387_ _2377_ _2388_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4435_ _1348_ _0944_ _0881_ _0859_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__3435__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4366_ _1362_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4892__A2 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6105_ mod.pc_1\[0\] _2827_ _2812_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3695__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3317_ mod.registers.r11\[0\] _3166_ _3168_ mod.registers.r8\[0\] _3169_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _0701_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2740_ _2755_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4266__I _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4644__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6938_ _0098_ net209 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6869_ _0029_ net151 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5825__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3345__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4332__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5560__I _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__A3 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__B1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3989__A4 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5060__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4571__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4323__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4220_ _0593_ _0598_ _0841_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4874__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ mod.registers.r13\[12\] _0929_ _0910_ mod.registers.r8\[12\] _1149_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5470__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ mod.registers.r12\[10\] _0716_ _0574_ mod.registers.r8\[10\] _1080_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_270 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__B1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_281 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_292 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6379__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _1965_ _1966_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ _0289_ net121 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3935_ _0914_ _0921_ _0927_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _0220_ net53 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3866_ _0456_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5605_ _2462_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6888__D _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6585_ _0151_ net128 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5645__I _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3797_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4562__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _2404_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6572__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _2203_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6303__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _1413_ _1407_ _1414_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5398_ _2318_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4865__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3668__A3 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4349_ _0945_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__B1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _1947_ _1948_ _1920_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__B1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4305__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5290__I _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4069__B1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6335__B _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ mod.registers.r13\[4\] _0689_ _0577_ mod.registers.r11\[4\] _0718_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3595__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__B2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ mod.pc_2\[10\] _3203_ _0641_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6370_ _1826_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3582_ _3153_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _2204_ _2274_ _2276_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6497__S _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ mod.registers.r1\[10\] _2205_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _1198_ _1199_ _0943_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _2123_ _2158_ _2159_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3713__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__C _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4134_ _0649_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6064__A4 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4065_ mod.registers.r5\[11\] _0897_ _0907_ mod.registers.r4\[11\] _0909_ mod.registers.r8\[11\]
+ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4075__A3 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A2 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4967_ _1863_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6706_ _0272_ net131 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3918_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3586__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ _1893_ _1606_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6637_ _0203_ net56 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3849_ _0846_ _0828_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _0134_ net129 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5519_ _2362_ _2412_ _2414_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _3088_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6288__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__B2 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4299__B1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout120 net123 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout131 net135 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout142 net143 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout153 net154 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout164 net167 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout175 net180 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout186 net191 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout197 net198 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__I _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6212__B2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4526__B2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6279__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6279__B2 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4565__S _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout184_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A2 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6203__B2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _1816_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4752_ _1050_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4765__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ _0678_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _1159_ _1175_ _1197_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3708__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A4 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ mod.des.des_dout\[2\] net18 _3045_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ _3238_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _2098_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3565_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5923__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5304_ mod.registers.r2\[2\] _2263_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3740__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout97_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _2940_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3496_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5235_ _2197_ _2204_ _2206_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4150__C1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ mod.registers.r1\[1\] _2137_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ _1112_ _1113_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ _3190_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5245__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4048_ mod.pc_2\[2\] _0594_ _1044_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__6760__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5999_ _1880_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3559__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4756__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4220__A3 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3618__I _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4508__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3716__C1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3731__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__I _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5484__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3495__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__B1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4598__I1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__B _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3970__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5172__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6633__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3350_ _3200_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _3131_ _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _0663_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6783__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3789__A2 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4450__A3 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5853_ _2383_ _2626_ _2630_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5918__I _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4738__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _0608_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5784_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4202__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _1520_ _1726_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__I3 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _1172_ _1154_ _1403_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3961__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6405_ _3026_ _1828_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3617_ _0411_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4597_ _1539_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5653__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ mod.pc_1\[13\] _2848_ _2987_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3548_ mod.registers.r11\[12\] _0497_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4269__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6267_ _2941_ _2944_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ mod.funct7\[0\] _0476_ _0447_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _2154_ _1988_ _2168_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6198_ mod.des.des_dout\[12\] _2888_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ mod.ins_ldr_3 mod.valid_out3 net15 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_28_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3901__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5218__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3348__I _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3952__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4179__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5457__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__I _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout147_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5393__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ _0852_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3943__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4451_ _1409_ _1231_ _1237_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5473__I _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3402_ _3253_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4382_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ mod.pc_1\[6\] _2834_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ mod.registers.r13\[0\] _3172_ _3176_ mod.registers.r14\[0\] _3184_ _3185_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_98_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1976_ _2775_ _2000_ _2780_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_105_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ mod.des.des_counter\[0\] _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ mod.pc_2\[6\] _1969_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ mod.registers.r14\[14\] _2660_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _0045_ net175 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _2612_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ mod.registers.r11\[11\] _2572_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4718_ _1130_ _1639_ _1091_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3934__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5698_ mod.registers.r10\[0\] _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6479__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4649_ _1208_ _1435_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ mod.pc_1\[7\] _2973_ _2971_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4111__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A2 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3689__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3689__B2 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4102__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3456__A4 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6821__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ mod.registers.r5\[7\] _0896_ _0578_ mod.registers.r10\[7\] _0949_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6073__B _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3613__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__I _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4372__I _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _0236_ net53 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3882_ _3211_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5621_ _2384_ _2474_ _2478_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4169__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5366__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _2345_ _2432_ _2435_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4503_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ mod.registers.r5\[11\] _2378_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4434_ _1242_ _1259_ _1428_ _1430_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4365_ _1226_ _1271_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4341__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3316_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1289_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2733_ _2765_ _2767_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6937_ _0097_ net208 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6868_ _0028_ net151 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5357__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ mod.registers.r12\[14\] _2606_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6799_ _0362_ net155 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__B _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3626__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__B1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3361__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6844__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__B2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4568__S _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ mod.registers.r12\[12\] _0904_ _0924_ mod.registers.r2\[12\] _0915_ mod.registers.r11\[12\]
+ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4081_ mod.registers.r3\[10\] _0680_ _0686_ mod.registers.r10\[10\] _1079_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_260 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3834__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_271 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3834__B2 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_282 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_293 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4983_ _1926_ _1967_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6722_ _0288_ net132 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4795__C1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3934_ mod.registers.r13\[15\] _0929_ _0931_ mod.registers.r9\[15\] _0932_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3865_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6653_ _0219_ net52 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5926__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__I _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _2460_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4011__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _0792_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6584_ _0150_ net127 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6717__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _2387_ _2418_ _2423_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ _2373_ _2363_ _2374_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4417_ _1413_ _1414_ _1407_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5511__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _2158_ _2319_ _2325_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4348_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4279_ _1276_ _0735_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4078__B2 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5578__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4250__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4305__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4069__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__B2 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B2 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4136__B _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3595__A3 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__B _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3650_ _0642_ _0645_ _0646_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6070__C _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3581_ mod.registers.r11\[1\] _0577_ _0578_ mod.registers.r10\[1\] _0579_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ mod.registers.r2\[8\] _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _2220_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6541__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__I _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4202_ _0943_ _1198_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_69_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ mod.registers.r1\[3\] _2137_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6049__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _1125_ _1129_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4064_ mod.registers.r3\[11\] _0899_ _0894_ mod.registers.r10\[11\] _1062_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3807__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout42_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4232__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4966_ mod.pc0\[5\] _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6705_ _0271_ net42 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3917_ _3165_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3586__A3 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5656__I _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _3210_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ _0202_ net57 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3848_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3779_ mod.registers.r7\[5\] _0750_ _0751_ mod.registers.r5\[5\] _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6567_ _0133_ net129 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3743__B1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5518_ mod.registers.r6\[4\] _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6498_ _3093_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6288__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5449_ _2164_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4299__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3904__I _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__B2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net113 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout132 net135 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout154 net161 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout165 net167 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout176 net180 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout187 net189 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5799__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__C _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3814__I _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3498__C1 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout177_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4462__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4751_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5962__A1 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__A2 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4380__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ _0564_ _0683_ _0695_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4682_ _1195_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ _3047_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3633_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4517__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3564_ _3226_ _0450_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6352_ _1821_ _2851_ _2998_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _2144_ _2261_ _2265_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6283_ _2948_ _2954_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3495_ _0435_ _0424_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ mod.registers.r1\[8\] _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__B1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4150__C2 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ mod.registers.r4\[9\] _0907_ _0917_ mod.registers.r14\[9\] _1114_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ _1893_ _1679_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6905__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ _0819_ _0820_ _0821_ _0822_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_72_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _1759_ _1878_ _1888_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5953__A1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4756__A2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _3190_ _1928_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5386__I _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4223__C _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _0185_ net52 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3716__B1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3716__C2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3634__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6130__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4692__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3495__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6585__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3955__B1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3280_ mod.instr_2\[14\] _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4435__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _1851_ _2668_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ mod.registers.r13\[10\] _2627_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4803_ _0609_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5935__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5783_ _2584_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4734_ _1072_ _1501_ _1728_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4665_ _1208_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5934__I _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ _2104_ _2992_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3616_ _0608_ _0429_ mod.registers.r2\[11\] _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5163__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _1036_ _1043_ _1052_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _1138_ _2920_ _2988_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3547_ mod.registers.r2\[12\] _0485_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6112__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3478_ _3141_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ _1347_ _2943_ _2938_ mod.instr\[9\] _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4994__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _1990_ _2179_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6197_ mod.instr\[12\] _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5148_ _2126_ _1344_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5079_ _2054_ _2062_ _2063_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4426__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4729__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3629__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5154__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__B1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__A2 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4417__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__I3 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ _1419_ _1421_ _1432_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6342__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ _3227_ _3229_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4381_ _0735_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _2811_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3332_ _3177_ _3178_ _3179_ _3182_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2757_ _2771_ _2776_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ _0586_ _1991_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4959__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__B2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _2394_ _2659_ _2662_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6884_ _0044_ net176 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5908__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ _2358_ _2613_ _2619_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ _2515_ _2571_ _2575_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5384__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _1637_ _1659_ _1679_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5697_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4648_ _1638_ _1641_ _1645_ _1609_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _1466_ _0860_ _1500_ _1042_ _3216_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _2678_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6249_ _2930_ _2931_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4647__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3912__I _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5072__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3359__I _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__B1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__B1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3689__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4099__C1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4139__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6354__B _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5749__I _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3613__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A1 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _3217_ _0462_ _0858_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ mod.registers.r8\[10\] _2475_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ mod.registers.r7\[0\] _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _0865_ _3207_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5482_ _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _1241_ _1261_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4364_ _1234_ _0862_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6079__B1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _2669_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3315_ _3159_ _3160_ _3142_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _1290_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ mod.pc\[4\] _2766_ _2748_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout72_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _0096_ net211 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6796__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _0027_ net152 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5818_ _2523_ _2605_ _2608_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _0361_ net156 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _2557_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3907__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3540__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3540__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6158__C _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4096__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3843__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__A2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4859__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__B _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__B2 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6669__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _1075_ _1076_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5284__A1 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4087__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_250 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_261 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A2 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_272 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_283 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_294 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5036__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__I _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A2 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _1929_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _0287_ net44 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3933_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__B1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__C2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _0218_ net90 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5339__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ _0563_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4547__B1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _2359_ _2461_ _2467_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6583_ _0149_ net128 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ mod.pc_2\[4\] _3204_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4011__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3727__I _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__I _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ mod.registers.r6\[11\] _2419_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ mod.registers.r5\[7\] _2364_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ _1231_ _1237_ _1409_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5511__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ mod.registers.r4\[3\] _2321_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4347_ mod.valid2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _0853_ _0722_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5275__A1 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4078__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _2698_ _1877_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3411__B _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _0079_ net59 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4250__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4002__A2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6013__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3761__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4896__C _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3372__I mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4069__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__I _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__I0 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _3161_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ mod.des.des_dout\[31\] _2207_ _2217_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__I1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4201_ _1191_ _1180_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3504__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _1111_ _1121_ _1123_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5257__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4063_ mod.registers.r7\[11\] _0892_ _0919_ mod.registers.r15\[11\] _1061_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3807__A2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1852_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4232__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _0270_ net45 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _0696_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3440__B1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ _1873_ _1874_ _1890_ _1892_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6635_ _0201_ net56 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3847_ _0463_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6834__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6566_ _0132_ net130 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3778_ mod.registers.r12\[5\] _0502_ _0494_ mod.registers.r15\[5\] _0776_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3743__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ _2406_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6497_ mod.des.des_dout\[16\] net19 _3089_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5448_ _2359_ _2348_ _2360_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4299__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4288__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout100 net102 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _2249_ _2308_ _2312_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout133 net135 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5248__A1 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout166 net167 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout177 net179 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout188 net189 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3920__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5847__I _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3734__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3498__B1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3498__C2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__I _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4462__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5411__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3701_ _0696_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4681_ _1662_ _1666_ _1667_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3277__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ mod.des.des_dout\[1\] net17 _3045_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3632_ mod.pc_2\[11\] _0453_ _0620_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5714__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ mod.rd_3\[1\] _2852_ _2097_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5492__I _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3563_ mod.pc_2\[12\] _3215_ _0553_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ mod.registers.r2\[1\] _2263_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6282_ _0585_ _2950_ _2953_ mod.instr\[15\] _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3494_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _2136_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ mod.des.des_dout\[22\] _2125_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4150__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4115_ mod.registers.r7\[9\] _0892_ _0923_ mod.registers.r2\[9\] _0915_ mod.registers.r11\[9\]
+ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _2079_ _2080_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _0814_ _0815_ _0816_ _0817_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_37_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4453__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3661__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _2730_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5667__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4948_ _1870_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4879_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6618_ _0184_ net56 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3716__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6549_ _0115_ net139 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6130__A2 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__B1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__B2 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5920_ _2667_ _2672_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _2380_ _2626_ _2629_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6092__B _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5487__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4802_ _1791_ _1794_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4733_ _1670_ _1729_ _1730_ _1394_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4664_ _1638_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5699__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _1777_ _3034_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3615_ _0612_ _0421_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4595_ _1373_ _1586_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6360__A2 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6334_ mod.pc_1\[12\] _2982_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3546_ mod.pc_2\[13\] _3205_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _2934_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__I _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3477_ _0468_ _0469_ _0470_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4123__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2160_ _2188_ _2189_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6196_ _2890_ _2891_ _2892_ _2884_ _2893_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5147_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _2064_ _1978_ _1981_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4426__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _1024_ _3203_ _1025_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_53_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3401__A3 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3645__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6351__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4362__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6552__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4114__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__I _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ mod.instr_2\[11\] mod.instr_2\[10\] _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout202_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4380_ _1264_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ mod.registers.r15\[0\] _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2742_ _2743_ _2001_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__B _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _0890_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ mod.registers.r14\[13\] _2660_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _0043_ net176 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5834_ mod.registers.r13\[3\] _2615_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6030__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ mod.registers.r11\[10\] _2572_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5384__A3 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _1694_ _1697_ _1700_ _1703_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4592__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5696_ _2529_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6575__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _1205_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3465__I _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4578_ _1572_ _1433_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _2975_ _2969_ _2976_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3529_ mod.registers.r8\[14\] _0487_ _0504_ mod.registers.r12\[14\] _0527_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5680__I _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A1 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _1816_ _2924_ _2928_ mod.instr\[4\] _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _2683_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3622__A3 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__I mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6021__A1 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4583__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__B2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3375__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__B2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6088__A1 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4099__B1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__C2 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__A1 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3613__A3 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__A2 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout152_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _0870_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_43_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6598__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4501_ _1288_ _1497_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5481_ _2227_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4432_ _1381_ _1429_ _1394_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4877__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4363_ _1297_ _1299_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6102_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__B2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3314_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4294_ _1267_ _1046_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2723_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout65_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0095_ net211 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _0026_ net165 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ mod.registers.r12\[13\] _2606_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _0360_ net149 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__B1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5748_ _2497_ _2558_ _2564_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _2235_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__S _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3540__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5817__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3679__I0 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__A1 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6740__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4005__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6890__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3531__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5808__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_240 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_251 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_262 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_273 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_284 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_295 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6233__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4981_ _1968_ _1969_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_45_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _0286_ net44 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3932_ _0711_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__B2 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6651_ _0217_ net56 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5495__I _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5602_ mod.registers.r8\[3\] _2463_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4547__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4547__B2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _0148_ net128 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3794_ _0786_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5533_ _2384_ _2418_ _2422_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4415_ _1108_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5395_ _2149_ _2319_ _2324_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6613__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ _0880_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _1270_ _1272_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ mod.pc\[3\] _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3286__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__A1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3589__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6918_ _0078_ net92 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _0009_ net168 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3918__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3761__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4010__I0 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4710__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6463__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__I1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6204__I mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout115_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _1159_ _1175_ _1195_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__C1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3504__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ mod.des.des_dout\[24\] _2151_ _2153_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6786__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ _0676_ _1107_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4062_ mod.registers.r12\[11\] _0905_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ mod.pc\[5\] _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _0269_ net42 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ mod.registers.r7\[15\] _0893_ _0895_ mod.registers.r10\[15\] _0912_ _0913_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3738__I _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _0571_ _0592_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3440__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3440__B2 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6114__I _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3846_ _0706_ _0571_ _0592_ _0597_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6634_ _0200_ net57 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6565_ _0131_ net138 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3777_ mod.registers.r9\[5\] _0506_ _0512_ mod.registers.r3\[5\] _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5516_ _2404_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3743__A2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _3092_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5447_ mod.registers.r5\[3\] _2350_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ mod.registers.r3\[14\] _2309_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout101 net102 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout134 net135 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4329_ _0883_ _1267_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout145 net200 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout156 net160 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout167 net182 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout189 net190 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4931__A1 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4479__I _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3383__I mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3498__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5239__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ mod.instr_2\[5\] _0697_ _0595_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _1378_ _1672_ _1673_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3631_ _0622_ _0625_ _0626_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6350_ _1818_ _2851_ _2997_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3562_ _0554_ _0555_ _0556_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3725__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5301_ _2135_ _2261_ _2264_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _2918_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3493_ _3246_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3293__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ _2139_ _1874_ _2132_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_57_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ mod.registers.r13\[9\] _0928_ _0925_ mod.registers.r1\[9\] _1112_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _3188_ _1152_ _2068_ _3190_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ _1037_ _1042_ _0440_ _0562_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6109__I _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3661__B2 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2725_ _2729_ _2731_ _2732_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _1749_ _1938_ _1939_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4878_ _1864_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5166__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _0183_ net89 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _0812_ _0825_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3716__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _0114_ net137 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6479_ _3062_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4677__B1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3931__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3378__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3404__B2 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__B _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4132__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout182_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__CLK net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5632__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A3 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4672__I _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ mod.registers.r13\[9\] _2627_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4801_ _1795_ _1796_ _1797_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5396__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _1427_ _1542_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4663_ _1660_ _1252_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5699__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3614_ _0411_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6402_ _3002_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ _0482_ _1590_ _1591_ _1508_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3545_ _0537_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6333_ _2963_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6264_ _2941_ _2942_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout95_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3476_ mod.registers.r13\[3\] _3172_ _3176_ mod.registers.r14\[3\] _0473_ _0474_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ mod.registers.r1\[6\] _2166_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4123__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__A1 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2718_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _1883_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ mod.pc\[11\] _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5623__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ _0805_ _0806_ _0807_ _0809_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__B1 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5979_ net11 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3926__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4362__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4114__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6847__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__C _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4353__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _3141_ _3180_ _3181_ _3174_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6368__B _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3571__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0888_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3616__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4813__C2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5902_ _2389_ _2659_ _2661_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6882_ _0042_ net193 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5369__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ _2355_ _2613_ _2618_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6030__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _2513_ _2571_ _2574_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _1452_ _1434_ _1699_ _1420_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5695_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4646_ _1238_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_163_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5541__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1288_ _1273_ _0872_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5961__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6316_ mod.pc_1\[6\] _2973_ _2971_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ mod.registers.r9\[14\] _0507_ _0495_ mod.registers.r15\[14\] _0526_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6247_ _2915_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3459_ _3225_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5844__A2 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ mod.des.des_dout\[7\] _2876_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ net12 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5201__I _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__A3 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5532__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4099__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__B2 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout145_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3566__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _1477_ _1424_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3782__B1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5480_ _2384_ _2377_ _2385_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4431_ _1288_ _1274_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4598__S _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _1306_ _1314_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6098__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6079__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _2669_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3313_ _3159_ _3160_ _3133_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4293_ _0812_ _1287_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _2757_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _0094_ net207 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4798__C1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _0025_ net164 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__C1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ _2519_ _2605_ _2607_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__B2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6796_ _0359_ net187 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5747_ mod.registers.r11\[3\] _2560_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5762__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3773__B1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _2517_ _2510_ _2518_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4317__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _1626_ _1364_ _1422_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3679__I1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4256__B _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4253__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4005__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4005__B2 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3603__I1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3764__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__B1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5808__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3819__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_230 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4492__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_241 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_252 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_263 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_274 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_285 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_296 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6233__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _0768_ _1950_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5992__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _0216_ net57 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _3206_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5601_ _2356_ _2461_ _2466_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5744__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4547__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _0147_ net137 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3793_ _0787_ _0788_ _0789_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5532_ mod.registers.r6\[10\] _2419_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _2194_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3507__B1 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4414_ _1407_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5394_ mod.registers.r4\[2\] _2321_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0874_ _1338_ _1339_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4276_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6908__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4855__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2733_ _2747_ _2749_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6472__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3286__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _0077_ net96 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__A1 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3589__A3 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ _0008_ net175 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0342_ net146 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6511__S _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6535__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4010__I1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6526__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__I _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__B2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__B1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__C2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _1088_ _1090_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6376__B _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__A2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4061_ _1034_ _1053_ _1054_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5009__A3 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4624__B _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5965__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _1947_ _1948_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0268_ net42 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3914_ _0901_ _0906_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4894_ _3187_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3440__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _0199_ net89 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3845_ _0842_ _0440_ _0826_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6564_ _0130_ net134 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ _0770_ _0771_ _0772_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5515_ _2359_ _2405_ _2411_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6517__I0 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ mod.des.des_dout\[15\] net18 _3089_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4940__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5446_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _2244_ _2308_ _2311_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout102 net108 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout135 net136 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4328_ _0853_ _0531_ _0451_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout146 net147 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout157 net160 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout168 net171 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout179 net180 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _1208_ _1255_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6880__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__S _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3498__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4695__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3670__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3630_ mod.registers.r1\[11\] _0510_ _0627_ mod.registers.r13\[11\] _0628_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6753__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _0557_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3574__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ mod.registers.r2\[0\] _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6124__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6280_ _2948_ _2952_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5231_ mod.des.des_dout\[29\] _2151_ _2200_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4686__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5162_ _1038_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ _0661_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5093_ _2075_ _2078_ _1870_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4438__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4044_ _3223_ _0844_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3661__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5938__A1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3749__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5995_ _2718_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6125__I _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ mod.pc\[4\] _1865_ _1867_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4610__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _3211_ _1581_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6616_ _0182_ net94 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ _0562_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6547_ _0113_ net137 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3484__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3759_ mod.registers.r6\[6\] _0604_ _0605_ mod.registers.r14\[6\] _0757_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6478_ _2386_ _3076_ _3081_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__B2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__I _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6626__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__B _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3404__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__I0 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A3 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5114__I _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout175_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _1769_ _1787_ _1785_ _1770_ _1788_ _1771_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _2316_ _2583_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4731_ _1309_ _1320_ _1283_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5784__I _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4662_ _1173_ _1159_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5148__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2684_ _3033_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3613_ _0420_ _0607_ mod.registers.r4\[11\] _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4593_ _1552_ _1435_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2985_ _2920_ _2986_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3544_ _0538_ _0539_ _0540_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6263_ _1348_ _2935_ _2938_ mod.instr\[8\] _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3475_ _0471_ _3178_ _3179_ _3182_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4659__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6194_ mod.des.des_dout\[11\] _2888_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4123__A3 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout88_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3882__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5076_ mod.pc0\[11\] _1958_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5959__I _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ _0800_ _0801_ _0802_ _0803_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_25_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _2685_ _2066_ _2717_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _1895_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4812__B _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5075__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__I mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3389__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4722__B _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4338__B1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4889__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3852__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3313__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6384__B _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__A1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6950_ _0110_ net201 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3616__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5901_ mod.registers.r14\[12\] _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _0041_ net183 mod.rd_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ mod.registers.r13\[2\] _2615_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ mod.registers.r11\[9\] _2572_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4041__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ _1709_ _1710_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5694_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4645_ _1239_ _1243_ _1642_ _1249_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _1340_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5541__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _1968_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4858__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _0522_ _0523_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6246_ _2922_ _2929_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3458_ mod.pc_2\[0\] _0453_ _0454_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _2674_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3389_ mod.instr_2\[13\] _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _2103_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__B1 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _1926_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4032__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__B2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3543__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__I0 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3543__B2 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__B1 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4271__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6424__S _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4452__B _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3782__A1 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3782__B2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _1359_ _1424_ _1426_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3534__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _1296_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6100_ _2818_ _2752_ _2821_ _2822_ _2823_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3312_ mod.registers.r10\[0\] _3161_ _3163_ mod.registers.r9\[0\] _3164_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4292_ _1035_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5287__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2761_ _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3298__B1 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__B1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6933_ _0093_ net209 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__B1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _0024_ net164 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__B1 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__C2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ mod.registers.r12\[12\] _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _0358_ net155 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _2495_ _2558_ _2563_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5762__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3773__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__B2 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ mod.registers.r9\[11\] _2511_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _1390_ _1267_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5514__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3525__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__B2 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4559_ _1317_ _1312_ _1272_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3492__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5278__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6229_ _2916_ _2856_ _2917_ _2858_ _2915_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6509__S _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3679__I2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4005__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__A1 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3603__I2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__B2 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__B2 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4713__B1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3819__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_220 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_231 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_242 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4492__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_253 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_264 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_275 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_286 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_297 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4244__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _3172_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _0850_ _3213_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3577__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5600_ mod.registers.r8\[2\] _2463_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6580_ _0146_ net133 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5744__A2 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3792_ mod.registers.r6\[4\] _3244_ _0750_ mod.registers.r7\[4\] _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ _2381_ _2418_ _2421_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ _2370_ _2363_ _2371_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3507__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3507__B2 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4413_ _1408_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5393_ _2144_ _2319_ _2323_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4180__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _0847_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6014_ mod.pc\[2\] _2737_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout70_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4483__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4235__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _0076_ net91 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5983__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3589__A4 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5188__B _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3487__I _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6847_ _0007_ net170 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _0341_ net146 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3746__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5729_ _2519_ _2550_ _2552_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6535__I1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4474__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A1 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3598__S _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4781__I mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6526__I1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6151__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5117__I _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4162__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__B2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _1055_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6682__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__B1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A2 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__I _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _1926_ _1949_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3913_ mod.registers.r4\[15\] _0908_ _0910_ mod.registers.r8\[15\] _0911_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6701_ _0267_ net68 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3976__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ _3126_ _1881_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6632_ _0198_ net95 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3844_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6563_ _0129_ net138 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3775_ mod.registers.r4\[5\] _3259_ _3220_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6390__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5514_ mod.registers.r6\[3\] _2407_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6517__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6494_ _3091_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5445_ _2157_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5376_ mod.registers.r3\[13\] _2309_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout103 net107 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6059__S _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout114 net124 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3770__I mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout125 net144 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout136 net142 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout158 net159 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4258_ _1194_ _1254_ _0942_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout169 net171 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ mod.registers.r11\[14\] _0916_ _0918_ mod.registers.r14\[14\] _1187_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5697__I _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6522__S _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5708__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3719__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3719__B2 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__I _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6555__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A2 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4695__A2 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5892__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3680__I _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3655__B1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__B _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__I0 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3670__A3 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__B2 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3855__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout120_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__I _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ mod.registers.r1\[12\] _0511_ _0490_ mod.registers.r13\[12\] _0558_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _0432_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4135__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _2171_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6387__B _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5883__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _1743_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _1108_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5092_ _2076_ _1876_ _1877_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4438__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _1038_ _0453_ _1039_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_37_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5938__A2 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ mod.pc\[0\] _2730_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3949__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4945_ mod.pc0\[4\] _1854_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4610__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6578__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3827_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6615_ _0181_ net94 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6141__I _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6546_ _0112_ net140 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3758_ mod.registers.r8\[6\] _3234_ _0602_ mod.registers.r10\[6\] _0756_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ mod.registers.r15\[11\] _3077_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5980__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ mod.registers.r10\[2\] _0686_ _0575_ mod.registers.r9\[2\] _0687_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4126__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _2134_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5874__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _2188_ _2296_ _2300_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6517__S _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3637__B1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4601__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4365__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__I1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__I _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5617__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__S _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3628__B1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3479__I0 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5093__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout168_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6720__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__B1 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4730_ _1630_ _1727_ _1073_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _1646_ _1657_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6345__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3585__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _1769_ _3028_ _3029_ _3015_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6870__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3612_ _0608_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _1588_ _1497_ _1589_ _1282_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ mod.pc_1\[11\] _2982_ _2979_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3543_ mod.registers.r7\[13\] _0516_ _0518_ mod.registers.r5\[13\] _0541_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4108__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3474_ mod.registers.r15\[3\] _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5213_ mod.des.des_dout\[27\] _2178_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _2674_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5144_ _2105_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5075_ _2040_ _2061_ _1966_ _1965_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ mod.pc_2\[3\] _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _2690_ mod.pc0\[11\] _2710_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _1749_ _1920_ _1921_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4812__C _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _0865_ _1349_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6336__A2 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A2 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _3111_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4320__S _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4338__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5838__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6263__B2 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3616__A3 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4813__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _2641_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ _0040_ net184 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6015__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _2352_ _2613_ _2617_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4577__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ _2509_ _2571_ _2573_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4713_ _1233_ _1630_ _1261_ _1236_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2258_ _2458_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1231_ _1237_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _1572_ _0452_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6616__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3526_ mod.registers.r1\[14\] _0511_ _0508_ mod.registers.r10\[14\] mod.registers.r14\[14\]
+ _0492_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6314_ _0769_ _2969_ _2974_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5829__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _1817_ _2924_ _2928_ mod.instr\[3\] _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3457_ _0416_ _0419_ _0427_ _0438_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5035__I mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ mod.instr\[7\] _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6766__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3388_ mod.registers.r8\[0\] _3234_ _3239_ mod.registers.r10\[0\] _3240_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _2104_ _2105_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _2041_ _2044_ _2042_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _0696_ _1001_ _1002_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4591__I1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3543__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A3 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4559__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6440__S _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3782__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout200_I mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1353_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3534__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6789__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _3158_ _3162_ _3145_ _3147_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1285_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _2742_ _2743_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5287__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3298__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5039__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6236__B2 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _0092_ net207 mod.des.des_dout\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__I0 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _0023_ net165 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__B2 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _2587_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6794_ _0357_ net156 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ mod.registers.r11\[2\] _2560_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4970__A1 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5676_ _2227_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4627_ _0812_ _1287_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3525__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _1304_ _1554_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _1464_ _1469_ _1222_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6475__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ mod.des.des_dout\[20\] _2866_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3679__I3 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6159_ mod.instr\[3\] _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6324__I _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__I3 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6931__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4013__I0 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_221 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_232 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_243 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_254 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_265 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_276 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_287 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_298 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A3 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout150_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3860_ _0704_ _0734_ _0849_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3791_ mod.registers.r13\[4\] _0433_ _0512_ mod.registers.r3\[4\] _0789_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ mod.registers.r6\[9\] _2419_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ mod.registers.r5\[6\] _2364_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _1022_ _1059_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3507__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4704__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ mod.registers.r4\[1\] _2321_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4274_ _0939_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _2695_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout63_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6915_ _0075_ net96 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3443__A1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _0409_ net175 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _0340_ net146 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3989_ _0885_ _0697_ mod.registers.r4\[6\] _0581_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3746__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ mod.registers.r10\[12\] _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5659_ _2187_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4171__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__I _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3985__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4302__I _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4162__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout198_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3673__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3673__B2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5414__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__B _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4961_ _1929_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _0266_ net69 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3912_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4892_ _1882_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6631_ _0197_ net90 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3843_ _0830_ _0463_ _0835_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6562_ _0128_ net134 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3774_ mod.registers.r2\[5\] _0483_ _3254_ mod.registers.r11\[5\] _0772_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5513_ _2356_ _2405_ _2410_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6493_ mod.des.des_dout\[14\] net17 _3089_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5308__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5444_ _2356_ _2348_ _2357_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5350__A1 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _2236_ _2308_ _2310_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout104 net107 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4326_ _0829_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout115 net119 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout137 net139 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout148 net149 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5102__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _0942_ _1194_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xfanout159 net160 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4188_ mod.registers.r12\[14\] _0905_ _0900_ mod.registers.r3\[14\] _0910_ mod.registers.r8\[14\]
+ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_27_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _0392_ net172 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5892__A2 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3655__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__B1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3490_ mod.registers.r2\[15\] _0485_ _0487_ mod.registers.r8\[15\] _0488_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__A1 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4135__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4967__I _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3871__I _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _1743_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5883__A2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ _1094_ _1107_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ mod.pc\[12\] _1866_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _0836_ _0837_ _0838_ _0839_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ _2723_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4207__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__A2 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1926_ _1928_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A3 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ mod.des.des_counter\[0\] _3120_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6614_ _0180_ net95 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _0813_ _3222_ _0818_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5571__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6545_ _0111_ _0003_ net206 mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3757_ _0740_ _3225_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_118_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _2383_ _3076_ _3080_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3688_ _3161_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5427_ _2255_ _2338_ _2343_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4126__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5874__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5358_ mod.registers.r3\[6\] _2297_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3885__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4309_ _0795_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5289_ mod.des.des_dout\[36\] _2178_ _2251_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3637__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3637__B2 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6533__S _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4365__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6672__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__I _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5865__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5617__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3628__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3628__B2 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3479__I1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__B1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ _1342_ _1641_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3611_ _3237_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5553__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _1211_ _1142_ _1135_ _1132_ _0796_ _0797_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _2057_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3542_ mod.registers.r1\[13\] _0511_ _0490_ mod.registers.r13\[13\] _0540_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5305__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4108__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3473_ mod.registers.r12\[3\] _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _2665_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _2180_ _2182_ _2184_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ mod.instr\[11\] _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5074_ _2056_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4025_ _0701_ _0825_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6417__I _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6545__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _2705_ _2050_ _2716_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4044__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4595__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ mod.pc\[3\] _1865_ _1748_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3398__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6152__I mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4858_ net13 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5544__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3809_ mod.registers.r9\[3\] _0422_ _0425_ mod.registers.r3\[3\] _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4789_ _3133_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6528_ net19 mod.des.des_dout\[29\] _3107_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _3062_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3858__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__S _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3686__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A2 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__S _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3313__A3 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout180_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3616__A4 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5830_ mod.registers.r13\[1\] _2615_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5774__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ mod.registers.r11\[8\] _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3596__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4712_ _1311_ _1375_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3785__B1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5692_ _2527_ _2520_ _2528_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1238_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_163_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ _1037_ _1042_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ mod.pc_1\[5\] _2973_ _2971_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3525_ mod.registers.r6\[14\] _0501_ _0497_ mod.registers.r11\[14\] _0523_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5829__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout93_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3456_ _3240_ _3248_ _3256_ _3263_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3304__A3 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ _2875_ _2867_ _2877_ _2872_ _2869_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3387_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5126_ mod.rd_3\[3\] _2100_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _2041_ _2042_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _1003_ _1004_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_84_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5765__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _2690_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__B1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6190__A1 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4740__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__I2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__A2 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4733__C _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4559__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6520__I _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3310_ mod.instr_2\[16\] _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _1286_ _1287_ _0452_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6484__A2 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3298__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__B _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6931_ _0091_ net210 mod.des.des_dout\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__I1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _0022_ net183 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5813_ _2585_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5747__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6793_ _0356_ net149 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3758__B1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5744_ _2493_ _2558_ _2562_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _2515_ _2510_ _2516_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4626_ _1509_ _1623_ _1264_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6733__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__B1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4557_ _1304_ _1326_ _1321_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3508_ _0422_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4488_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6227_ mod.instr\[20\] _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6475__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3439_ _3177_ _0434_ _0435_ _0436_ _3183_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6158_ _2862_ _2675_ _2864_ _2859_ _2823_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _2052_ _1694_ _1697_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4238__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ _1980_ _2074_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6541__S _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4013__I1 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 net30 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6466__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_222 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6218__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_233 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_244 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_255 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_266 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_277 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_288 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_299 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6606__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3452__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3790_ mod.registers.r8\[4\] _0486_ _0747_ mod.registers.r1\[4\] _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6756__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6154__B2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4411_ _1110_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4165__B1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2135_ _2319_ _2322_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _3192_ _3207_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6457__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4273_ _0458_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6012_ _2740_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

