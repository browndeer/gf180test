// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire net91;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net92;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net93;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net129;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net130;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net131;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net159;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net160;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net161;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net162;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net163;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net164;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire \mod.clk ;
 wire \mod.des.des_counter[0] ;
 wire \mod.des.des_counter[1] ;
 wire \mod.des.des_counter[2] ;
 wire \mod.des.des_din[24] ;
 wire \mod.des.des_dout[0] ;
 wire \mod.des.des_dout[10] ;
 wire \mod.des.des_dout[11] ;
 wire \mod.des.des_dout[12] ;
 wire \mod.des.des_dout[13] ;
 wire \mod.des.des_dout[14] ;
 wire \mod.des.des_dout[15] ;
 wire \mod.des.des_dout[16] ;
 wire \mod.des.des_dout[17] ;
 wire \mod.des.des_dout[18] ;
 wire \mod.des.des_dout[19] ;
 wire \mod.des.des_dout[1] ;
 wire \mod.des.des_dout[20] ;
 wire \mod.des.des_dout[21] ;
 wire \mod.des.des_dout[22] ;
 wire \mod.des.des_dout[23] ;
 wire \mod.des.des_dout[2] ;
 wire \mod.des.des_dout[3] ;
 wire \mod.des.des_dout[4] ;
 wire \mod.des.des_dout[5] ;
 wire \mod.des.des_dout[6] ;
 wire \mod.des.des_dout[7] ;
 wire \mod.des.des_dout[8] ;
 wire \mod.des.des_dout[9] ;
 wire \mod.funct3[0] ;
 wire \mod.funct3[1] ;
 wire \mod.funct3[2] ;
 wire \mod.ins_ldr_3 ;
 wire \mod.instr[0] ;
 wire \mod.instr[10] ;
 wire \mod.instr[11] ;
 wire \mod.instr[12] ;
 wire \mod.instr[13] ;
 wire \mod.instr[14] ;
 wire \mod.instr[15] ;
 wire \mod.instr[1] ;
 wire \mod.instr[2] ;
 wire \mod.instr[3] ;
 wire \mod.instr[4] ;
 wire \mod.instr[5] ;
 wire \mod.instr[6] ;
 wire \mod.instr[7] ;
 wire \mod.instr[8] ;
 wire \mod.instr[9] ;
 wire \mod.instr_2[0] ;
 wire \mod.instr_2[10] ;
 wire \mod.instr_2[11] ;
 wire \mod.instr_2[12] ;
 wire \mod.instr_2[13] ;
 wire \mod.instr_2[14] ;
 wire \mod.instr_2[15] ;
 wire \mod.instr_2[1] ;
 wire \mod.instr_2[2] ;
 wire \mod.instr_2[3] ;
 wire \mod.instr_2[4] ;
 wire \mod.instr_2[5] ;
 wire \mod.instr_2[9] ;
 wire \mod.ldr_hzd[0] ;
 wire \mod.ldr_hzd[1] ;
 wire \mod.ldr_hzd[2] ;
 wire \mod.ldr_hzd[3] ;
 wire \mod.ldr_hzd[4] ;
 wire \mod.ldr_hzd[5] ;
 wire \mod.ldr_hzd[6] ;
 wire \mod.ldr_hzd[7] ;
 wire \mod.pc0[0] ;
 wire \mod.pc0[1] ;
 wire \mod.pc0[2] ;
 wire \mod.pc0[3] ;
 wire \mod.pc0[4] ;
 wire \mod.pc0[5] ;
 wire \mod.pc[0] ;
 wire \mod.pc[1] ;
 wire \mod.pc[2] ;
 wire \mod.pc[3] ;
 wire \mod.pc[4] ;
 wire \mod.pc[5] ;
 wire \mod.pc_1[0] ;
 wire \mod.pc_1[1] ;
 wire \mod.pc_1[2] ;
 wire \mod.pc_1[3] ;
 wire \mod.pc_1[4] ;
 wire \mod.pc_1[5] ;
 wire \mod.pc_2[0] ;
 wire \mod.pc_2[1] ;
 wire \mod.pc_2[2] ;
 wire \mod.pc_2[3] ;
 wire \mod.pc_2[4] ;
 wire \mod.pc_2[5] ;
 wire \mod.rd_3[0] ;
 wire \mod.rd_3[1] ;
 wire \mod.rd_3[2] ;
 wire \mod.registers.r1[0] ;
 wire \mod.registers.r1[1] ;
 wire \mod.registers.r1[2] ;
 wire \mod.registers.r1[3] ;
 wire \mod.registers.r1[4] ;
 wire \mod.registers.r1[5] ;
 wire \mod.registers.r1[6] ;
 wire \mod.registers.r1[7] ;
 wire \mod.registers.r2[0] ;
 wire \mod.registers.r2[1] ;
 wire \mod.registers.r2[2] ;
 wire \mod.registers.r2[3] ;
 wire \mod.registers.r2[4] ;
 wire \mod.registers.r2[5] ;
 wire \mod.registers.r2[6] ;
 wire \mod.registers.r2[7] ;
 wire \mod.registers.r3[0] ;
 wire \mod.registers.r3[1] ;
 wire \mod.registers.r3[2] ;
 wire \mod.registers.r3[3] ;
 wire \mod.registers.r3[4] ;
 wire \mod.registers.r3[5] ;
 wire \mod.registers.r3[6] ;
 wire \mod.registers.r3[7] ;
 wire \mod.registers.r4[0] ;
 wire \mod.registers.r4[1] ;
 wire \mod.registers.r4[2] ;
 wire \mod.registers.r4[3] ;
 wire \mod.registers.r4[4] ;
 wire \mod.registers.r4[5] ;
 wire \mod.registers.r4[6] ;
 wire \mod.registers.r4[7] ;
 wire \mod.registers.r5[0] ;
 wire \mod.registers.r5[1] ;
 wire \mod.registers.r5[2] ;
 wire \mod.registers.r5[3] ;
 wire \mod.registers.r5[4] ;
 wire \mod.registers.r5[5] ;
 wire \mod.registers.r5[6] ;
 wire \mod.registers.r5[7] ;
 wire \mod.registers.r6[0] ;
 wire \mod.registers.r6[1] ;
 wire \mod.registers.r6[2] ;
 wire \mod.registers.r6[3] ;
 wire \mod.registers.r6[4] ;
 wire \mod.registers.r6[5] ;
 wire \mod.registers.r6[6] ;
 wire \mod.registers.r6[7] ;
 wire \mod.registers.r7[0] ;
 wire \mod.registers.r7[1] ;
 wire \mod.registers.r7[2] ;
 wire \mod.registers.r7[3] ;
 wire \mod.registers.r7[4] ;
 wire \mod.registers.r7[5] ;
 wire \mod.registers.r7[6] ;
 wire \mod.registers.r7[7] ;
 wire \mod.ri_3 ;
 wire \mod.valid0 ;
 wire \mod.valid1 ;
 wire \mod.valid2 ;
 wire \mod.valid_out3 ;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1176_ (.I(\mod.des.des_counter[1] ),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1177_ (.A1(\mod.des.des_counter[0] ),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1178_ (.A1(net26),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1179_ (.I(_0527_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1180_ (.I(\mod.des.des_counter[0] ),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1181_ (.I(_0528_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1182_ (.I(\mod.des.des_counter[0] ),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1183_ (.I(\mod.des.des_counter[1] ),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1184_ (.A1(_0529_),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1185_ (.A1(_0528_),
    .A2(_0525_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1186_ (.I(_0532_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1187_ (.A1(_0531_),
    .A2(_0533_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1188_ (.I(\mod.des.des_counter[2] ),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1189_ (.A1(_0534_),
    .A2(_0526_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1190_ (.I(_0535_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1191_ (.A1(_0529_),
    .A2(_0525_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1192_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1193_ (.I(\mod.valid2 ),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1194_ (.I(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1195_ (.I(\mod.funct3[1] ),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1196_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1197_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1198_ (.I(\mod.funct3[0] ),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1199_ (.I(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1200_ (.I(\mod.instr_2[15] ),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1201_ (.I(\mod.instr_2[2] ),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1202_ (.I(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1203_ (.I(\mod.instr_2[0] ),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1204_ (.I(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1205_ (.I(\mod.instr_2[1] ),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1206_ (.A1(_0547_),
    .A2(_0549_),
    .B(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1207_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1208_ (.A1(_0545_),
    .A2(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1209_ (.I(_0552_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1210_ (.I(\mod.instr_2[13] ),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1211_ (.I(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1212_ (.I(\mod.instr_2[12] ),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1213_ (.A1(_0556_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1214_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1215_ (.I(\mod.instr_2[12] ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1216_ (.A1(\mod.instr_2[13] ),
    .A2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1217_ (.I(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1218_ (.A1(_0555_),
    .A2(_0557_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1219_ (.I(_0563_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1220_ (.A1(\mod.registers.r2[6] ),
    .A2(_0559_),
    .B1(_0562_),
    .B2(\mod.registers.r1[6] ),
    .C1(_0564_),
    .C2(\mod.registers.r3[6] ),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1221_ (.A1(_0554_),
    .A2(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1222_ (.A1(_0553_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1223_ (.I(\mod.instr_2[11] ),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1224_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1225_ (.I(\mod.instr_2[10] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1226_ (.I(\mod.instr_2[9] ),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1227_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1228_ (.I(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1229_ (.I(_0570_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1230_ (.A1(\mod.instr_2[11] ),
    .A2(_0574_),
    .A3(_0571_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1231_ (.I(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1232_ (.I(\mod.instr_2[11] ),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1233_ (.I(\mod.instr_2[10] ),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1234_ (.A1(_0577_),
    .A2(_0578_),
    .A3(_0571_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1235_ (.I(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1236_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1237_ (.A1(\mod.registers.r7[6] ),
    .A2(_0573_),
    .B1(_0576_),
    .B2(\mod.registers.r3[6] ),
    .C1(_0581_),
    .C2(\mod.registers.r1[6] ),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1238_ (.A1(_0568_),
    .A2(_0578_),
    .A3(_0571_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1239_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1240_ (.I(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1241_ (.I(\mod.instr_2[9] ),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1242_ (.A1(_0569_),
    .A2(_0574_),
    .A3(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1243_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1244_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1245_ (.A1(\mod.registers.r5[6] ),
    .A2(_0585_),
    .B1(_0589_),
    .B2(\mod.registers.r6[6] ),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1246_ (.A1(\mod.instr_2[11] ),
    .A2(_0574_),
    .A3(_0586_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1247_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1248_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1249_ (.A1(_0569_),
    .A2(_0578_),
    .A3(_0586_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1250_ (.I(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1251_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1252_ (.A1(\mod.registers.r2[6] ),
    .A2(_0593_),
    .B1(_0596_),
    .B2(\mod.registers.r4[6] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1253_ (.A1(_0582_),
    .A2(_0590_),
    .A3(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1254_ (.A1(_0567_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1255_ (.A1(_0567_),
    .A2(_0598_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1256_ (.A1(_0599_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1257_ (.A1(\mod.registers.r2[5] ),
    .A2(_0559_),
    .B1(_0562_),
    .B2(\mod.registers.r1[5] ),
    .C1(_0564_),
    .C2(\mod.registers.r3[5] ),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1258_ (.I(_0551_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1259_ (.A1(\mod.instr_2[15] ),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1260_ (.A1(_0554_),
    .A2(_0602_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1261_ (.I(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1262_ (.A1(\mod.registers.r3[5] ),
    .A2(_0576_),
    .B1(_0585_),
    .B2(\mod.registers.r5[5] ),
    .C1(\mod.registers.r6[5] ),
    .C2(_0589_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1263_ (.A1(\mod.registers.r7[5] ),
    .A2(_0573_),
    .B1(_0581_),
    .B2(\mod.registers.r1[5] ),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1264_ (.A1(\mod.registers.r2[5] ),
    .A2(_0593_),
    .B1(_0596_),
    .B2(\mod.registers.r4[5] ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1265_ (.A1(_0607_),
    .A2(_0608_),
    .A3(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1266_ (.I(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1267_ (.A1(_0606_),
    .A2(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1268_ (.A1(\mod.registers.r2[4] ),
    .A2(_0558_),
    .B1(_0562_),
    .B2(\mod.registers.r1[4] ),
    .C1(_0563_),
    .C2(\mod.registers.r3[4] ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1269_ (.A1(_0603_),
    .A2(_0613_),
    .B(_0604_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1270_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1271_ (.I(_0575_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1272_ (.A1(\mod.registers.r7[4] ),
    .A2(_0573_),
    .B1(_0585_),
    .B2(\mod.registers.r5[4] ),
    .C1(_0616_),
    .C2(\mod.registers.r3[4] ),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1273_ (.A1(\mod.registers.r2[4] ),
    .A2(_0593_),
    .B1(_0596_),
    .B2(\mod.registers.r4[4] ),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1274_ (.A1(\mod.registers.r1[4] ),
    .A2(_0581_),
    .B1(_0589_),
    .B2(\mod.registers.r6[4] ),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1275_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1276_ (.I(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1277_ (.A1(_0615_),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1278_ (.A1(_0614_),
    .A2(_0621_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1279_ (.A1(_0622_),
    .A2(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1280_ (.I(_0572_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1281_ (.A1(\mod.registers.r7[3] ),
    .A2(_0625_),
    .B1(_0580_),
    .B2(\mod.registers.r1[3] ),
    .C1(_0588_),
    .C2(\mod.registers.r6[3] ),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1282_ (.A1(\mod.registers.r3[3] ),
    .A2(_0616_),
    .B1(_0595_),
    .B2(\mod.registers.r4[3] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1283_ (.A1(\mod.registers.r5[3] ),
    .A2(_0584_),
    .B1(_0592_),
    .B2(\mod.registers.r2[3] ),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1284_ (.A1(_0626_),
    .A2(_0627_),
    .A3(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1285_ (.I(_0546_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1286_ (.I(_0548_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1287_ (.I(\mod.instr_2[1] ),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1288_ (.A1(_0630_),
    .A2(_0631_),
    .B(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1289_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1290_ (.I(_0586_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1291_ (.A1(_0546_),
    .A2(_0548_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1292_ (.A1(\mod.funct3[2] ),
    .A2(\mod.instr_2[1] ),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1293_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1294_ (.A1(_0636_),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1295_ (.I0(\mod.instr_2[14] ),
    .I1(_0635_),
    .S(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1296_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1297_ (.A1(_0546_),
    .A2(\mod.instr_2[0] ),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1298_ (.A1(\mod.instr_2[1] ),
    .A2(_0641_),
    .B1(_0642_),
    .B2(_0637_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1299_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1300_ (.I0(_0640_),
    .I1(\mod.instr_2[15] ),
    .S(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1301_ (.A1(\mod.registers.r2[3] ),
    .A2(_0558_),
    .B1(_0561_),
    .B2(\mod.registers.r1[3] ),
    .C1(_0563_),
    .C2(\mod.registers.r3[3] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1302_ (.A1(_0633_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1303_ (.A1(_0634_),
    .A2(_0645_),
    .B(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1304_ (.A1(_0629_),
    .A2(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1305_ (.A1(\mod.registers.r3[2] ),
    .A2(_0616_),
    .B1(_0595_),
    .B2(\mod.registers.r4[2] ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1306_ (.A1(\mod.registers.r5[2] ),
    .A2(_0584_),
    .B1(_0592_),
    .B2(\mod.registers.r2[2] ),
    .C1(_0588_),
    .C2(\mod.registers.r6[2] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1307_ (.A1(\mod.registers.r7[2] ),
    .A2(_0625_),
    .B1(_0580_),
    .B2(\mod.registers.r1[2] ),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1308_ (.A1(_0650_),
    .A2(_0651_),
    .A3(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1309_ (.I(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1310_ (.I(\mod.instr_2[5] ),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1311_ (.A1(\mod.funct3[2] ),
    .A2(_0632_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1312_ (.A1(_0630_),
    .A2(_0548_),
    .B(\mod.funct3[2] ),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1313_ (.A1(_0655_),
    .A2(_0642_),
    .A3(_0656_),
    .B(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1314_ (.I0(_0658_),
    .I1(\mod.instr_2[14] ),
    .S(_0643_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1315_ (.I(\mod.instr_2[13] ),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1316_ (.I(_0560_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1317_ (.A1(_0660_),
    .A2(_0661_),
    .A3(\mod.registers.r2[2] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1318_ (.A1(\mod.registers.r3[2] ),
    .A2(_0563_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1319_ (.A1(_0556_),
    .A2(_0557_),
    .A3(\mod.registers.r1[2] ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1320_ (.A1(_0662_),
    .A2(_0663_),
    .A3(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1321_ (.I0(_0659_),
    .I1(_0665_),
    .S(_0551_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1322_ (.I(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1323_ (.A1(_0654_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1324_ (.A1(\mod.registers.r2[1] ),
    .A2(_0591_),
    .B1(_0594_),
    .B2(\mod.registers.r4[1] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1325_ (.A1(\mod.registers.r1[1] ),
    .A2(_0579_),
    .B1(_0583_),
    .B2(\mod.registers.r5[1] ),
    .C1(\mod.registers.r6[1] ),
    .C2(_0587_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1326_ (.A1(\mod.registers.r7[1] ),
    .A2(_0625_),
    .B1(_0616_),
    .B2(\mod.registers.r3[1] ),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1327_ (.A1(_0669_),
    .A2(_0670_),
    .A3(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1328_ (.I(_0636_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1329_ (.A1(\mod.instr_2[4] ),
    .A2(_0673_),
    .A3(_0638_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1330_ (.A1(\mod.funct3[1] ),
    .A2(_0639_),
    .B(_0674_),
    .C(_0643_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1331_ (.A1(_0556_),
    .A2(_0644_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1332_ (.A1(_0660_),
    .A2(_0560_),
    .A3(\mod.registers.r2[1] ),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1333_ (.I(\mod.registers.r1[1] ),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1334_ (.A1(_0555_),
    .A2(_0557_),
    .A3(\mod.registers.r3[1] ),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1335_ (.A1(_0660_),
    .A2(_0560_),
    .A3(_0678_),
    .B(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1336_ (.A1(_0677_),
    .A2(_0680_),
    .B(_0551_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1337_ (.A1(_0603_),
    .A2(_0675_),
    .A3(_0676_),
    .B(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1338_ (.A1(_0672_),
    .A2(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1339_ (.A1(\mod.registers.r3[0] ),
    .A2(_0576_),
    .B1(_0595_),
    .B2(\mod.registers.r4[0] ),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1340_ (.A1(\mod.registers.r5[0] ),
    .A2(_0584_),
    .B1(_0588_),
    .B2(\mod.registers.r6[0] ),
    .C1(\mod.registers.r2[0] ),
    .C2(_0592_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1341_ (.A1(\mod.registers.r7[0] ),
    .A2(_0625_),
    .B1(_0580_),
    .B2(\mod.registers.r1[0] ),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1342_ (.A1(_0684_),
    .A2(_0685_),
    .A3(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1343_ (.I(\mod.instr_2[3] ),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1344_ (.I(_0642_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1345_ (.A1(_0688_),
    .A2(_0689_),
    .A3(_0656_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1346_ (.A1(\mod.funct3[0] ),
    .A2(_0639_),
    .B(_0690_),
    .C(_0644_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1347_ (.A1(_0661_),
    .A2(_0644_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1348_ (.I(_0555_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1349_ (.A1(_0693_),
    .A2(_0661_),
    .A3(\mod.registers.r2[0] ),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1350_ (.I(\mod.registers.r1[0] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1351_ (.I(\mod.instr_2[12] ),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1352_ (.A1(_0660_),
    .A2(_0696_),
    .A3(\mod.registers.r3[0] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1353_ (.A1(_0693_),
    .A2(_0661_),
    .A3(_0695_),
    .B(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1354_ (.A1(_0694_),
    .A2(_0698_),
    .B(_0603_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1355_ (.A1(_0552_),
    .A2(_0691_),
    .A3(_0692_),
    .B(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1356_ (.A1(_0687_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1357_ (.A1(_0672_),
    .A2(_0682_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1358_ (.A1(_0653_),
    .A2(_0666_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1359_ (.A1(_0683_),
    .A2(_0701_),
    .B(_0702_),
    .C(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1360_ (.I(_0629_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1361_ (.I(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1362_ (.I(_0648_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1363_ (.A1(_0706_),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1364_ (.A1(_0649_),
    .A2(_0668_),
    .A3(_0704_),
    .B(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1365_ (.A1(_0615_),
    .A2(_0620_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1366_ (.I(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1367_ (.A1(_0606_),
    .A2(_0611_),
    .B1(_0624_),
    .B2(_0709_),
    .C(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1368_ (.I(_0554_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1369_ (.A1(_0713_),
    .A2(_0565_),
    .B(_0604_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1370_ (.A1(_0601_),
    .A2(_0612_),
    .A3(_0712_),
    .B1(_0598_),
    .B2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1371_ (.A1(\mod.registers.r2[7] ),
    .A2(_0559_),
    .B1(_0562_),
    .B2(\mod.registers.r1[7] ),
    .C1(_0564_),
    .C2(\mod.registers.r3[7] ),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1372_ (.A1(_0554_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1373_ (.A1(_0553_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1374_ (.A1(\mod.registers.r7[7] ),
    .A2(_0573_),
    .B1(_0576_),
    .B2(\mod.registers.r3[7] ),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1375_ (.A1(\mod.registers.r1[7] ),
    .A2(_0581_),
    .B1(_0585_),
    .B2(\mod.registers.r5[7] ),
    .C1(\mod.registers.r6[7] ),
    .C2(_0589_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1376_ (.A1(\mod.registers.r2[7] ),
    .A2(_0593_),
    .B1(_0596_),
    .B2(\mod.registers.r4[7] ),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1377_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1378_ (.A1(_0718_),
    .A2(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1379_ (.I(_0722_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1380_ (.A1(_0553_),
    .A2(_0717_),
    .A3(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1381_ (.A1(_0715_),
    .A2(_0723_),
    .B(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1382_ (.A1(_0544_),
    .A2(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1383_ (.A1(_0542_),
    .A2(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1384_ (.I(\mod.funct3[2] ),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1385_ (.I(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1386_ (.I(_0544_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1387_ (.A1(_0715_),
    .A2(_0723_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1388_ (.A1(_0599_),
    .A2(_0600_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1389_ (.A1(_0612_),
    .A2(_0712_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1390_ (.A1(_0733_),
    .A2(_0612_),
    .A3(_0712_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1391_ (.A1(_0606_),
    .A2(_0610_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1392_ (.A1(_0605_),
    .A2(_0611_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1393_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1394_ (.A1(_0624_),
    .A2(_0709_),
    .B(_0711_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1395_ (.A1(_0738_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1396_ (.I(_0624_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1397_ (.A1(_0741_),
    .A2(_0709_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1398_ (.I(_0649_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1399_ (.I(_0683_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1400_ (.I(_0687_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1401_ (.I(_0552_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1402_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1403_ (.A1(_0694_),
    .A2(_0698_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1404_ (.A1(_0746_),
    .A2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1405_ (.A1(_0746_),
    .A2(_0747_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1406_ (.A1(_0745_),
    .A2(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1407_ (.I(_0750_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1408_ (.A1(_0745_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1409_ (.A1(_0751_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1410_ (.A1(_0703_),
    .A2(_0668_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1411_ (.A1(_0743_),
    .A2(_0744_),
    .A3(_0754_),
    .A4(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1412_ (.A1(_0742_),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1413_ (.A1(_0734_),
    .A2(_0735_),
    .A3(_0740_),
    .A4(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1414_ (.I(_0541_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1415_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1416_ (.A1(_0731_),
    .A2(_0732_),
    .A3(_0758_),
    .B(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1417_ (.A1(_0730_),
    .A2(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1418_ (.I(\mod.funct3[0] ),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1419_ (.I(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1420_ (.I(_0723_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1421_ (.A1(_0715_),
    .A2(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1422_ (.A1(_0764_),
    .A2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1423_ (.I(_0732_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1424_ (.I(_0729_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1425_ (.A1(_0731_),
    .A2(_0768_),
    .B(_0769_),
    .C(_0760_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1426_ (.A1(_0729_),
    .A2(_0541_),
    .A3(_0763_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1427_ (.A1(_0768_),
    .A2(_0758_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1428_ (.A1(_0632_),
    .A2(_0673_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1429_ (.I(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1430_ (.A1(_0767_),
    .A2(_0770_),
    .B(_0772_),
    .C(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1431_ (.I(_0630_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1432_ (.A1(_0776_),
    .A2(_0549_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1433_ (.A1(_0728_),
    .A2(_0762_),
    .A3(_0775_),
    .B(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(_0539_),
    .A2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1435_ (.I(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1436_ (.I(\mod.pc[0] ),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1437_ (.I(\mod.ldr_hzd[0] ),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1438_ (.I(_0635_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1439_ (.I(\mod.ldr_hzd[1] ),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1440_ (.A1(_0784_),
    .A2(_0783_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1441_ (.A1(_0782_),
    .A2(_0783_),
    .B(_0785_),
    .C(_0574_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1442_ (.I(_0578_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1443_ (.I(\mod.ldr_hzd[3] ),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1444_ (.A1(\mod.ldr_hzd[2] ),
    .A2(_0635_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1445_ (.A1(_0788_),
    .A2(_0783_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1446_ (.A1(_0787_),
    .A2(_0790_),
    .B(_0577_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1447_ (.I0(\mod.ldr_hzd[4] ),
    .I1(\mod.ldr_hzd[5] ),
    .I2(\mod.ldr_hzd[6] ),
    .I3(\mod.ldr_hzd[7] ),
    .S0(_0635_),
    .S1(_0787_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1448_ (.A1(_0569_),
    .A2(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1449_ (.A1(_0786_),
    .A2(_0791_),
    .B(_0776_),
    .C(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(\mod.ldr_hzd[2] ),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1451_ (.A1(\mod.ldr_hzd[0] ),
    .A2(_0696_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1452_ (.A1(_0784_),
    .A2(_0696_),
    .B(_0796_),
    .C(_0693_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1453_ (.A1(_0795_),
    .A2(_0559_),
    .B1(_0564_),
    .B2(\mod.ldr_hzd[3] ),
    .C(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1454_ (.A1(_0630_),
    .A2(_0549_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1455_ (.I(_0632_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1456_ (.A1(_0776_),
    .A2(_0800_),
    .A3(_0631_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1457_ (.A1(_0777_),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1458_ (.A1(_0799_),
    .A2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1459_ (.A1(_0689_),
    .A2(_0638_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(\mod.instr_2[3] ),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1461_ (.I(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1462_ (.A1(_0788_),
    .A2(_0805_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1463_ (.I(\mod.instr_2[4] ),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1464_ (.A1(_0795_),
    .A2(_0806_),
    .B(_0807_),
    .C(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1465_ (.A1(\mod.instr_2[4] ),
    .A2(_0688_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1466_ (.A1(\mod.instr_2[4] ),
    .A2(_0805_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1467_ (.A1(\mod.ldr_hzd[1] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(_0782_),
    .C(\mod.instr_2[5] ),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1468_ (.I(_0688_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1469_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_0805_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1470_ (.A1(\mod.ldr_hzd[7] ),
    .A2(_0813_),
    .B(_0814_),
    .C(_0808_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1471_ (.A1(\mod.ldr_hzd[5] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(\mod.ldr_hzd[4] ),
    .C(_0655_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1472_ (.A1(_0809_),
    .A2(_0812_),
    .B1(_0815_),
    .B2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1473_ (.A1(_0804_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1474_ (.A1(_0639_),
    .A2(_0798_),
    .B(_0803_),
    .C(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1475_ (.A1(\mod.ldr_hzd[3] ),
    .A2(_0795_),
    .A3(\mod.ldr_hzd[1] ),
    .A4(_0782_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1476_ (.A1(\mod.ldr_hzd[7] ),
    .A2(\mod.ldr_hzd[6] ),
    .A3(\mod.ldr_hzd[5] ),
    .A4(\mod.ldr_hzd[4] ),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1477_ (.A1(_0820_),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1478_ (.A1(_0794_),
    .A2(_0819_),
    .B(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1479_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1480_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1482_ (.A1(\mod.pc0[0] ),
    .A2(_0825_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1483_ (.A1(_0781_),
    .A2(_0826_),
    .B(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1484_ (.A1(_0800_),
    .A2(_0777_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1485_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1486_ (.I0(_0768_),
    .I1(_0726_),
    .S(_0763_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1487_ (.I(_0673_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1488_ (.I(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1489_ (.A1(_0769_),
    .A2(_0760_),
    .A3(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1490_ (.I(_0707_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1491_ (.I(_0667_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1492_ (.I(_0700_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1493_ (.I(_0615_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1494_ (.A1(_0598_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1495_ (.A1(_0837_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1496_ (.I(_0615_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1497_ (.I(_0750_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1498_ (.A1(_0841_),
    .A2(_0842_),
    .A3(_0722_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1499_ (.A1(_0840_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1500_ (.I(_0700_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1501_ (.A1(_0845_),
    .A2(_0710_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1502_ (.A1(_0610_),
    .A2(_0838_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1503_ (.A1(_0842_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1504_ (.A1(_0846_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1505_ (.A1(_0675_),
    .A2(_0676_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1506_ (.A1(_0677_),
    .A2(_0680_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1507_ (.A1(_0746_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1508_ (.A1(_0746_),
    .A2(_0850_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1509_ (.I(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1510_ (.I0(_0844_),
    .I1(_0849_),
    .S(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1511_ (.A1(_0836_),
    .A2(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1512_ (.I(_0845_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1513_ (.A1(_0838_),
    .A2(_0654_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1514_ (.A1(_0857_),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1515_ (.I(_0752_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1516_ (.A1(_0838_),
    .A2(_0705_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1517_ (.A1(_0860_),
    .A2(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1518_ (.A1(_0859_),
    .A2(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1519_ (.I(_0672_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1520_ (.A1(_0841_),
    .A2(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1521_ (.A1(_0860_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1522_ (.A1(_0854_),
    .A2(_0866_),
    .B(_0836_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1523_ (.A1(_0841_),
    .A2(_0745_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1524_ (.I(_0682_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1525_ (.A1(_0869_),
    .A2(_0837_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1526_ (.A1(_0868_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1527_ (.A1(_0854_),
    .A2(_0863_),
    .B(_0867_),
    .C(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_0730_),
    .A2(_0673_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1529_ (.A1(_0763_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1530_ (.A1(_0541_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1531_ (.A1(_0835_),
    .A2(_0856_),
    .A3(_0872_),
    .A4(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1532_ (.A1(_0634_),
    .A2(_0659_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1533_ (.A1(_0713_),
    .A2(_0665_),
    .B(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1534_ (.A1(_0729_),
    .A2(_0540_),
    .A3(_0832_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1535_ (.A1(_0543_),
    .A2(_0707_),
    .A3(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1536_ (.I(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1537_ (.A1(_0878_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1538_ (.A1(_0871_),
    .A2(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1539_ (.A1(_0540_),
    .A2(_0873_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1540_ (.A1(_0540_),
    .A2(_0543_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1541_ (.A1(_0832_),
    .A2(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1542_ (.A1(_0543_),
    .A2(_0884_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(_0753_),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1544_ (.A1(_0751_),
    .A2(_0884_),
    .B1(_0886_),
    .B2(_0754_),
    .C(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1545_ (.A1(_0883_),
    .A2(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1546_ (.A1(_0876_),
    .A2(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1547_ (.A1(_0831_),
    .A2(_0834_),
    .B(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1548_ (.I(\mod.pc_2[0] ),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1549_ (.A1(_0691_),
    .A2(_0692_),
    .B(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1550_ (.A1(\mod.pc_2[0] ),
    .A2(_0747_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1551_ (.A1(_0894_),
    .A2(_0895_),
    .B(_0829_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1552_ (.A1(_0830_),
    .A2(_0892_),
    .B(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1553_ (.A1(_0538_),
    .A2(_0778_),
    .A3(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1554_ (.A1(_0780_),
    .A2(_0828_),
    .B(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1555_ (.I(_0525_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1556_ (.A1(_0000_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1557_ (.I(_0873_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1558_ (.A1(_0902_),
    .A2(_0886_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1559_ (.I(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1560_ (.A1(_0744_),
    .A2(_0701_),
    .B(_0702_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1561_ (.A1(_0864_),
    .A2(_0853_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1562_ (.A1(_0864_),
    .A2(_0853_),
    .B(_0745_),
    .C(_0750_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1563_ (.A1(_0906_),
    .A2(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1564_ (.A1(_0545_),
    .A2(_0799_),
    .A3(_0638_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1565_ (.A1(_0773_),
    .A2(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1566_ (.I0(_0905_),
    .I1(_0908_),
    .S(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1567_ (.A1(_0755_),
    .A2(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1568_ (.A1(_0860_),
    .A2(_0868_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1569_ (.A1(_0859_),
    .A2(_0866_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1570_ (.I(_0854_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1571_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1572_ (.I0(_0913_),
    .I1(_0914_),
    .S(_0916_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1573_ (.A1(_0882_),
    .A2(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1574_ (.I(_0875_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1575_ (.A1(_0724_),
    .A2(_0910_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1576_ (.A1(_0836_),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1577_ (.I(_0835_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1578_ (.A1(_0667_),
    .A2(_0853_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1579_ (.A1(_0667_),
    .A2(_0869_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1580_ (.A1(_0840_),
    .A2(_0843_),
    .B(_0915_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1581_ (.I(_0836_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1582_ (.A1(_0849_),
    .A2(_0923_),
    .B1(_0924_),
    .B2(_0863_),
    .C1(_0925_),
    .C2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1583_ (.A1(_0922_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1584_ (.A1(_0916_),
    .A2(_0921_),
    .B(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1585_ (.A1(_0902_),
    .A2(_0885_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1586_ (.A1(_0759_),
    .A2(_0874_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1587_ (.A1(_0654_),
    .A2(_0878_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1588_ (.A1(_0654_),
    .A2(_0878_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1589_ (.A1(_0931_),
    .A2(_0932_),
    .B1(_0933_),
    .B2(_0887_),
    .C(_0903_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1590_ (.A1(_0755_),
    .A2(_0930_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1591_ (.A1(_0919_),
    .A2(_0929_),
    .B(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1592_ (.A1(_0904_),
    .A2(_0912_),
    .B1(_0918_),
    .B2(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_0901_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1594_ (.I(\mod.des.des_din[24] ),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1595_ (.A1(_0939_),
    .A2(_0530_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1596_ (.A1(_0532_),
    .A2(_0665_),
    .B1(_0940_),
    .B2(_0000_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1597_ (.A1(_0537_),
    .A2(_0899_),
    .B1(_0938_),
    .B2(_0941_),
    .ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1598_ (.I(\mod.valid2 ),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1599_ (.A1(_0732_),
    .A2(_0758_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1600_ (.A1(_0731_),
    .A2(_0768_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1601_ (.A1(_0764_),
    .A2(_0766_),
    .B(_0730_),
    .C(_0542_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1602_ (.A1(_0943_),
    .A2(_0771_),
    .B1(_0944_),
    .B2(_0945_),
    .C(_0773_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1603_ (.A1(_0542_),
    .A2(_0727_),
    .B1(_0761_),
    .B2(_0730_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1604_ (.A1(_0547_),
    .A2(_0631_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1605_ (.A1(_0946_),
    .A2(_0947_),
    .B(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1606_ (.A1(_0942_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1607_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1608_ (.I0(\mod.pc0[1] ),
    .I1(\mod.pc[1] ),
    .S(_0825_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1609_ (.I(\mod.pc_2[1] ),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1610_ (.I(_0850_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1611_ (.A1(_0953_),
    .A2(_0954_),
    .A3(_0895_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1612_ (.I(_0869_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1613_ (.A1(_0956_),
    .A2(_0857_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1614_ (.I(_0878_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1615_ (.A1(_0752_),
    .A2(_0839_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1616_ (.A1(_0845_),
    .A2(_0847_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1617_ (.A1(_0959_),
    .A2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1618_ (.A1(_0841_),
    .A2(_0845_),
    .A3(_0722_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1619_ (.A1(_0869_),
    .A2(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1620_ (.A1(_0956_),
    .A2(_0961_),
    .B(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1621_ (.A1(_0752_),
    .A2(_0861_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1622_ (.A1(_0842_),
    .A2(_0711_),
    .B(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(_0842_),
    .A2(_0865_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1624_ (.A1(_0837_),
    .A2(_0858_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1625_ (.A1(_0967_),
    .A2(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1626_ (.A1(_0923_),
    .A2(_0966_),
    .B1(_0969_),
    .B2(_0924_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1627_ (.A1(_0958_),
    .A2(_0964_),
    .B(_0970_),
    .C(_0835_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1628_ (.A1(_0921_),
    .A2(_0957_),
    .B(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1629_ (.A1(_0875_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(_0860_),
    .A2(_0868_),
    .B(_0967_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1631_ (.A1(_0956_),
    .A2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1632_ (.A1(_0958_),
    .A2(_0881_),
    .A3(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1633_ (.A1(_0864_),
    .A2(_0915_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1634_ (.A1(_0744_),
    .A2(_0930_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1635_ (.A1(_0977_),
    .A2(_0887_),
    .B1(_0931_),
    .B2(_0906_),
    .C(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1636_ (.A1(_0837_),
    .A2(_0910_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1637_ (.A1(_0744_),
    .A2(_0701_),
    .A3(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1638_ (.A1(_0903_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1639_ (.A1(_0973_),
    .A2(_0976_),
    .A3(_0979_),
    .A4(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1640_ (.I0(_0955_),
    .I1(_0983_),
    .S(_0830_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1641_ (.A1(_0538_),
    .A2(_0778_),
    .A3(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1642_ (.A1(_0951_),
    .A2(_0952_),
    .B(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1643_ (.I(_0923_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1644_ (.A1(_0915_),
    .A2(_0962_),
    .B(_0958_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1645_ (.A1(_0987_),
    .A2(_0961_),
    .B1(_0966_),
    .B2(_0924_),
    .C(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1646_ (.A1(_0922_),
    .A2(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1647_ (.A1(_0870_),
    .A2(_0921_),
    .B(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(_0919_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1649_ (.I(_0657_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1650_ (.A1(_0649_),
    .A2(_0993_),
    .B1(_0885_),
    .B2(_0833_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1651_ (.I(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1652_ (.I(_0764_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1653_ (.A1(_0705_),
    .A2(_0707_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1654_ (.A1(_0705_),
    .A2(_0835_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1655_ (.A1(_0996_),
    .A2(_0997_),
    .B(_0884_),
    .C(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1656_ (.A1(_0965_),
    .A2(_0968_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1657_ (.I0(_0974_),
    .I1(_1000_),
    .S(_0916_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1658_ (.A1(_0882_),
    .A2(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1659_ (.A1(_0995_),
    .A2(_0999_),
    .A3(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1660_ (.I(_0910_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1661_ (.A1(_0908_),
    .A2(_0932_),
    .B(_0933_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1662_ (.A1(_0668_),
    .A2(_0704_),
    .A3(_1004_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1663_ (.A1(_1004_),
    .A2(_1005_),
    .B(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1664_ (.A1(_0743_),
    .A2(_1007_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1665_ (.A1(_0992_),
    .A2(_1003_),
    .B1(_1008_),
    .B2(_0904_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1666_ (.I(_0529_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1667_ (.A1(_1010_),
    .A2(_0646_),
    .B(_0900_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1668_ (.A1(_0000_),
    .A2(_1009_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1669_ (.A1(_0537_),
    .A2(_0986_),
    .B(_1012_),
    .ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1670_ (.I(\mod.pc[2] ),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1671_ (.I(_0824_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1672_ (.A1(\mod.pc0[2] ),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1673_ (.A1(_1013_),
    .A2(_0826_),
    .B(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1674_ (.I(_0779_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1675_ (.I(_0830_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1676_ (.I(\mod.pc_2[2] ),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1677_ (.I(_0659_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1678_ (.A1(\mod.pc_2[1] ),
    .A2(_0954_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1679_ (.A1(_0953_),
    .A2(_0954_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1680_ (.A1(_0895_),
    .A2(_1021_),
    .B(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1681_ (.A1(_1019_),
    .A2(_1020_),
    .A3(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1682_ (.A1(_1018_),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1683_ (.A1(_1018_),
    .A2(_0937_),
    .B(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1684_ (.A1(_1017_),
    .A2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1685_ (.A1(_0780_),
    .A2(_1016_),
    .B(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1686_ (.A1(_0528_),
    .A2(_0530_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1687_ (.I(_1004_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1688_ (.A1(_0997_),
    .A2(_1005_),
    .B(_0998_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(_0773_),
    .A2(_0909_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1690_ (.A1(_0741_),
    .A2(_1031_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1691_ (.A1(_0741_),
    .A2(_1031_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1692_ (.A1(_0742_),
    .A2(_1030_),
    .B(_0904_),
    .C(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1693_ (.I(_0958_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1694_ (.A1(_0922_),
    .A2(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1695_ (.A1(_0855_),
    .A2(_1037_),
    .B(_0921_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1696_ (.I(_0924_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1697_ (.A1(_0846_),
    .A2(_0862_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1699_ (.A1(_0926_),
    .A2(_0871_),
    .B1(_0987_),
    .B2(_0914_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1700_ (.A1(_0881_),
    .A2(_1041_),
    .A3(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1701_ (.I(_0622_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1702_ (.A1(_1044_),
    .A2(_0887_),
    .B1(_0931_),
    .B2(_0623_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1703_ (.A1(_0741_),
    .A2(_0930_),
    .B(_1043_),
    .C(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1704_ (.A1(_0919_),
    .A2(_1038_),
    .B(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1705_ (.A1(_1035_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1706_ (.A1(_0901_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1707_ (.A1(_0533_),
    .A2(_0613_),
    .B1(_1028_),
    .B2(_1029_),
    .C(_1049_),
    .ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1708_ (.I(_0830_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1709_ (.I(\mod.pc_2[3] ),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1710_ (.I(_0645_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1711_ (.A1(_1019_),
    .A2(_1020_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1712_ (.A1(\mod.pc_2[2] ),
    .A2(_1020_),
    .B(_1023_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1713_ (.A1(_1053_),
    .A2(_1054_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1714_ (.A1(_1051_),
    .A2(_1052_),
    .A3(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1715_ (.A1(_1018_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1716_ (.A1(_1050_),
    .A2(_1009_),
    .B(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1717_ (.I0(\mod.pc0[3] ),
    .I1(\mod.pc[3] ),
    .S(_0824_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1718_ (.I(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1719_ (.I0(_1058_),
    .I1(_1060_),
    .S(_1017_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1720_ (.A1(_0740_),
    .A2(_1030_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1721_ (.A1(_0623_),
    .A2(_1031_),
    .B(_1044_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1722_ (.A1(_0738_),
    .A2(_1063_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1723_ (.A1(_1032_),
    .A2(_1064_),
    .B(_0904_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1724_ (.A1(_0760_),
    .A2(_0996_),
    .A3(_0902_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1725_ (.A1(_0922_),
    .A2(_1036_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1726_ (.A1(_1036_),
    .A2(_0957_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1727_ (.A1(_1067_),
    .A2(_0964_),
    .B1(_1068_),
    .B2(_0920_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1728_ (.A1(_1066_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1729_ (.A1(_0993_),
    .A2(_0738_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1730_ (.I(_0542_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1731_ (.I(_0736_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1732_ (.A1(_0996_),
    .A2(_0737_),
    .B(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1733_ (.A1(_1072_),
    .A2(_0902_),
    .A3(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1734_ (.A1(_0857_),
    .A2(_0711_),
    .B(_0960_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1735_ (.A1(_0956_),
    .A2(_1000_),
    .B1(_1076_),
    .B2(_1039_),
    .C(_0880_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1736_ (.A1(_1036_),
    .A2(_0975_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1737_ (.A1(_0886_),
    .A2(_1071_),
    .B(_1075_),
    .C(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1738_ (.A1(_1062_),
    .A2(_1065_),
    .B1(_1070_),
    .B2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1739_ (.A1(_0529_),
    .A2(_0602_),
    .B(_0900_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1740_ (.I(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1741_ (.A1(_0536_),
    .A2(_1061_),
    .B1(_1080_),
    .B2(_1010_),
    .C(_1082_),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1742_ (.I(\mod.pc[4] ),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1743_ (.A1(\mod.pc0[4] ),
    .A2(_1014_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1744_ (.A1(_1083_),
    .A2(_0826_),
    .B(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1745_ (.A1(_0689_),
    .A2(_0713_),
    .B(_0545_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1746_ (.A1(_0787_),
    .A2(_0832_),
    .A3(_0634_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1747_ (.A1(_1086_),
    .A2(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1748_ (.A1(\mod.pc_2[4] ),
    .A2(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1749_ (.A1(\mod.pc_2[3] ),
    .A2(_1052_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(_1051_),
    .A2(_1052_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1751_ (.A1(_1090_),
    .A2(_1055_),
    .B(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(_1089_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1753_ (.A1(_1089_),
    .A2(_1092_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1754_ (.A1(_1018_),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1755_ (.A1(_1050_),
    .A2(_1048_),
    .B1(_1093_),
    .B2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1756_ (.A1(_1017_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1757_ (.A1(_0780_),
    .A2(_1085_),
    .B(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1758_ (.A1(_1073_),
    .A2(_1063_),
    .B(_0737_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1759_ (.A1(_1073_),
    .A2(_1063_),
    .B(_0737_),
    .C(_0733_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1760_ (.A1(_1032_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1761_ (.A1(_0601_),
    .A2(_1099_),
    .B(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1762_ (.A1(_0734_),
    .A2(_0735_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_0833_),
    .A2(_0771_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1764_ (.A1(_1103_),
    .A2(_1032_),
    .B(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1765_ (.A1(_0724_),
    .A2(_1039_),
    .A3(_1004_),
    .B1(_0925_),
    .B2(_1037_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1766_ (.I(_1039_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1767_ (.A1(_0987_),
    .A2(_1040_),
    .B(_0880_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1768_ (.A1(_0840_),
    .A2(_0848_),
    .A3(_1107_),
    .B(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1769_ (.A1(_0926_),
    .A2(_0917_),
    .B(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1770_ (.I(_0599_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1771_ (.A1(_0764_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1772_ (.A1(_1072_),
    .A2(_1111_),
    .B(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1773_ (.A1(_0600_),
    .A2(_0993_),
    .A3(_1113_),
    .B(_1104_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1774_ (.A1(_0919_),
    .A2(_1106_),
    .B(_1110_),
    .C(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1775_ (.A1(_1102_),
    .A2(_1105_),
    .B(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1776_ (.A1(_0901_),
    .A2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1777_ (.A1(_0533_),
    .A2(_0565_),
    .B1(_1098_),
    .B2(_1029_),
    .C(_1117_),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1778_ (.I(\mod.pc[5] ),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1779_ (.A1(\mod.pc0[5] ),
    .A2(_1014_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1780_ (.A1(_1118_),
    .A2(_0826_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(\mod.pc_2[4] ),
    .A2(_1088_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1782_ (.A1(_1121_),
    .A2(_1093_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1783_ (.A1(_0577_),
    .A2(_0833_),
    .A3(_0634_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1784_ (.A1(_1086_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1785_ (.A1(\mod.pc_2[5] ),
    .A2(_1122_),
    .A3(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1786_ (.A1(_1050_),
    .A2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1787_ (.A1(_1050_),
    .A2(_1080_),
    .B(_1126_),
    .C(_0779_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1788_ (.A1(_0780_),
    .A2(_1120_),
    .B(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1789_ (.A1(_0987_),
    .A2(_1076_),
    .B(_0880_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1790_ (.A1(_1107_),
    .A2(_0962_),
    .A3(_0959_),
    .B(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1791_ (.A1(_0926_),
    .A2(_1001_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1792_ (.A1(_0916_),
    .A2(_1067_),
    .A3(_0962_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1793_ (.A1(_0857_),
    .A2(_1107_),
    .B(_0920_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1794_ (.A1(_1132_),
    .A2(_1133_),
    .B(_1066_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1795_ (.A1(_0718_),
    .A2(_0724_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1796_ (.A1(_1072_),
    .A2(_1135_),
    .B1(_0765_),
    .B2(_0731_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1797_ (.A1(_0993_),
    .A2(_1136_),
    .B(_1104_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1798_ (.A1(_1111_),
    .A2(_1100_),
    .B(_0765_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1799_ (.A1(_1111_),
    .A2(_0765_),
    .A3(_1100_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1800_ (.A1(_1030_),
    .A2(_1138_),
    .A3(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1801_ (.A1(_0766_),
    .A2(_1030_),
    .B(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1802_ (.A1(_1131_),
    .A2(_1134_),
    .A3(_1137_),
    .B1(_1141_),
    .B2(_1104_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1803_ (.A1(_0531_),
    .A2(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1804_ (.A1(_0533_),
    .A2(_0716_),
    .B1(_1128_),
    .B2(_1029_),
    .C(_1143_),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1805_ (.A1(_0538_),
    .A2(_0823_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1806_ (.A1(_0800_),
    .A2(_0532_),
    .A3(_0689_),
    .A4(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1807_ (.A1(_1010_),
    .A2(_0748_),
    .B(_0900_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1808_ (.A1(_0769_),
    .A2(_1145_),
    .B(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1809_ (.A1(_0537_),
    .A2(_0892_),
    .B(_1147_),
    .ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1810_ (.A1(_1010_),
    .A2(_0851_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1811_ (.A1(_0530_),
    .A2(_1148_),
    .B(_1145_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1812_ (.A1(_0537_),
    .A2(_0983_),
    .B(_1149_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1813_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1814_ (.I(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1815_ (.I0(\mod.rd_3[1] ),
    .I1(_0808_),
    .S(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1816_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1817_ (.I(_1153_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(\mod.rd_3[0] ),
    .A2(_1153_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1819_ (.A1(_0813_),
    .A2(_1154_),
    .B(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1820_ (.I(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1821_ (.A1(_1152_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1822_ (.I(_0655_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1823_ (.I(_1150_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1824_ (.A1(\mod.rd_3[2] ),
    .A2(_1151_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1825_ (.A1(_0803_),
    .A2(_1144_),
    .B(_1150_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1826_ (.A1(net7),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1827_ (.A1(_1159_),
    .A2(_1160_),
    .B(_1161_),
    .C(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_1158_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1829_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1830_ (.I(_1154_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1831_ (.I(_0801_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1832_ (.I(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1833_ (.I(_0777_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1834_ (.I(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1835_ (.A1(_1171_),
    .A2(_1048_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1836_ (.I(_0948_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(\mod.pc_2[4] ),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1838_ (.A1(_1169_),
    .A2(_1172_),
    .A3(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1839_ (.A1(_0954_),
    .A2(_1169_),
    .B(_1160_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1840_ (.I(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1841_ (.A1(\mod.des.des_dout[20] ),
    .A2(_1167_),
    .B1(_1175_),
    .B2(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1842_ (.I(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1843_ (.I(_1165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1844_ (.A1(\mod.registers.r5[4] ),
    .A2(_0166_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1845_ (.A1(_1166_),
    .A2(_0165_),
    .B(_0167_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(\mod.des.des_dout[21] ),
    .A2(_1167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1847_ (.A1(\mod.pc_2[5] ),
    .A2(_0948_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1848_ (.A1(_1173_),
    .A2(_1080_),
    .B(_0169_),
    .C(_1168_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1849_ (.A1(_1020_),
    .A2(_1169_),
    .B(_1160_),
    .C(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_0168_),
    .A2(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1851_ (.I(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1852_ (.I(_1165_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1853_ (.I0(_0173_),
    .I1(\mod.registers.r5[5] ),
    .S(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1854_ (.I(_0175_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1855_ (.I(_1151_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1856_ (.I(_1052_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1857_ (.I(_1168_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1858_ (.A1(_1171_),
    .A2(_0178_),
    .A3(_1116_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1859_ (.A1(_0177_),
    .A2(_1169_),
    .B(_0176_),
    .C(_0179_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1860_ (.A1(\mod.des.des_dout[22] ),
    .A2(_0176_),
    .B(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1861_ (.I(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1862_ (.A1(\mod.registers.r5[6] ),
    .A2(_0166_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1863_ (.A1(_1166_),
    .A2(_0182_),
    .B(_0183_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1864_ (.A1(_0178_),
    .A2(_1086_),
    .A3(_1087_),
    .B1(_1142_),
    .B2(_0802_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1865_ (.I0(\mod.des.des_dout[23] ),
    .I1(_0184_),
    .S(_0176_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1866_ (.I(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1867_ (.I0(_0186_),
    .I1(\mod.registers.r5[7] ),
    .S(_0174_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1868_ (.I(_0187_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1869_ (.I(\mod.des.des_dout[16] ),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1870_ (.A1(_0178_),
    .A2(_1151_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1871_ (.I0(_0893_),
    .I1(_0892_),
    .S(_1170_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1872_ (.A1(_0188_),
    .A2(_0176_),
    .B1(_0189_),
    .B2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1873_ (.I(_0191_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1874_ (.I(_1152_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1875_ (.A1(_0193_),
    .A2(_1156_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1876_ (.A1(_1164_),
    .A2(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1877_ (.I(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1878_ (.I0(_0192_),
    .I1(\mod.registers.r6[0] ),
    .S(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1879_ (.I(_0197_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1880_ (.I(_0195_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1881_ (.A1(_0953_),
    .A2(_1170_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1882_ (.A1(_1171_),
    .A2(_0983_),
    .B(_0189_),
    .C(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1883_ (.A1(\mod.des.des_dout[17] ),
    .A2(_1167_),
    .B(_0200_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1884_ (.I(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1885_ (.I(_0195_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1886_ (.A1(\mod.registers.r6[1] ),
    .A2(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1887_ (.A1(_0198_),
    .A2(_0202_),
    .B(_0204_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1888_ (.A1(_1173_),
    .A2(_0937_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1889_ (.A1(_1019_),
    .A2(_1171_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1890_ (.A1(_0189_),
    .A2(_0205_),
    .A3(_0206_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1891_ (.A1(\mod.des.des_dout[18] ),
    .A2(_1167_),
    .B(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1892_ (.I(_0208_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1893_ (.A1(\mod.registers.r6[2] ),
    .A2(_0203_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1894_ (.A1(_0198_),
    .A2(_0209_),
    .B(_0210_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1895_ (.A1(_1173_),
    .A2(_1009_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1896_ (.A1(_1051_),
    .A2(_1170_),
    .B(_1168_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1897_ (.A1(_0691_),
    .A2(_0692_),
    .A3(_0178_),
    .B1(_0211_),
    .B2(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1898_ (.I0(\mod.des.des_dout[19] ),
    .I1(_0213_),
    .S(_1160_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1899_ (.I(_0214_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1900_ (.I0(_0215_),
    .I1(\mod.registers.r6[3] ),
    .S(_0196_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1901_ (.I(_0216_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1902_ (.A1(\mod.registers.r6[4] ),
    .A2(_0203_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1903_ (.A1(_0165_),
    .A2(_0198_),
    .B(_0217_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1904_ (.I0(_0173_),
    .I1(\mod.registers.r6[5] ),
    .S(_0196_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1905_ (.I(_0218_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1906_ (.A1(\mod.registers.r6[6] ),
    .A2(_0203_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1907_ (.A1(_0182_),
    .A2(_0198_),
    .B(_0219_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1908_ (.I0(_0186_),
    .I1(\mod.registers.r6[7] ),
    .S(_0196_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1909_ (.I(_0220_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1910_ (.I(net9),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1911_ (.I(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1912_ (.I(_0222_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1913_ (.I(net9),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1914_ (.I(_0223_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1915_ (.I(_0224_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1916_ (.I(_0225_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1917_ (.I(_0225_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1918_ (.I(net7),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1919_ (.A1(_0226_),
    .A2(_0825_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1920_ (.I(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1921_ (.A1(_0950_),
    .A2(_0823_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(\mod.valid0 ),
    .A2(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1923_ (.I(net9),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1924_ (.I(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1925_ (.A1(_0228_),
    .A2(_0230_),
    .B(_0232_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1926_ (.A1(_0534_),
    .A2(_0526_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1927_ (.I(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1928_ (.I0(\mod.des.des_dout[18] ),
    .I1(net1),
    .S(_0234_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1929_ (.I(_0235_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1930_ (.I0(\mod.des.des_dout[19] ),
    .I1(net2),
    .S(_0234_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1931_ (.I(_0236_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1932_ (.I0(\mod.des.des_dout[20] ),
    .I1(net3),
    .S(_0234_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(_0237_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1934_ (.I0(\mod.des.des_dout[21] ),
    .I1(net4),
    .S(_0234_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1935_ (.I(_0238_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1936_ (.I0(\mod.des.des_dout[22] ),
    .I1(net5),
    .S(_0233_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1937_ (.I(_0239_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1938_ (.I0(\mod.des.des_dout[23] ),
    .I1(net6),
    .S(_0233_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1939_ (.I(_0240_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1940_ (.A1(net7),
    .A2(_0823_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1941_ (.A1(\mod.valid0 ),
    .A2(_0241_),
    .A3(_0229_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1942_ (.I(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1943_ (.I(_0227_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1944_ (.A1(\mod.valid1 ),
    .A2(_0244_),
    .A3(_0229_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1945_ (.I(_0231_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1946_ (.A1(_0243_),
    .A2(_0245_),
    .B(_0246_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1947_ (.I(_0226_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1948_ (.I(_0247_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1949_ (.I(_0226_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1950_ (.I(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1951_ (.A1(_0250_),
    .A2(\mod.pc0[0] ),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1952_ (.I(_0231_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1953_ (.A1(_0248_),
    .A2(_0899_),
    .B(_0251_),
    .C(_0252_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1954_ (.A1(_0250_),
    .A2(\mod.pc0[1] ),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1955_ (.A1(_0248_),
    .A2(_0986_),
    .B(_0253_),
    .C(_0252_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1956_ (.I(_0249_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1957_ (.A1(_0254_),
    .A2(\mod.pc0[2] ),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1958_ (.A1(_0248_),
    .A2(_1028_),
    .B(_0255_),
    .C(_0252_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1959_ (.A1(_0254_),
    .A2(\mod.pc0[3] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1960_ (.I(_0231_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1961_ (.A1(_0248_),
    .A2(_1061_),
    .B(_0256_),
    .C(_0257_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1962_ (.A1(_0254_),
    .A2(\mod.pc0[4] ),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1963_ (.A1(_0250_),
    .A2(_1098_),
    .B(_0258_),
    .C(_0257_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1964_ (.A1(_0254_),
    .A2(\mod.pc0[5] ),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1965_ (.A1(_0250_),
    .A2(_1128_),
    .B(_0259_),
    .C(_0257_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1966_ (.A1(_0951_),
    .A2(_0824_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1967_ (.A1(_0226_),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1968_ (.I(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1969_ (.I(_0261_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1970_ (.A1(_0539_),
    .A2(_0778_),
    .B(_0781_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1971_ (.A1(_0898_),
    .A2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1972_ (.I(_0221_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1973_ (.I(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1974_ (.A1(_0263_),
    .A2(_0265_),
    .B(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1975_ (.A1(_0781_),
    .A2(_0262_),
    .B(_0268_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1976_ (.I(\mod.pc[1] ),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1977_ (.A1(_0942_),
    .A2(_0949_),
    .B(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1978_ (.A1(_0898_),
    .A2(_0264_),
    .B(_0985_),
    .C(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1979_ (.I(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1980_ (.A1(_0985_),
    .A2(_0270_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1981_ (.A1(_0265_),
    .A2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1982_ (.A1(_0272_),
    .A2(_0274_),
    .B(_0263_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1983_ (.A1(_0269_),
    .A2(_0262_),
    .B(_0275_),
    .C(_0257_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1984_ (.I0(_1013_),
    .I1(_1026_),
    .S(_0950_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1985_ (.A1(_0272_),
    .A2(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1986_ (.A1(_0271_),
    .A2(_0276_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1987_ (.A1(_0277_),
    .A2(_0278_),
    .B(_0263_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1988_ (.I(_0223_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1989_ (.A1(_1013_),
    .A2(_0262_),
    .B(_0279_),
    .C(_0280_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1990_ (.A1(_0249_),
    .A2(_0260_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1991_ (.I(\mod.pc[3] ),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1992_ (.I0(_0282_),
    .I1(_1058_),
    .S(_0951_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1993_ (.A1(_0278_),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(\mod.pc[3] ),
    .A2(_0281_),
    .B(_0267_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1995_ (.A1(_0281_),
    .A2(_0284_),
    .B(_0285_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1996_ (.A1(_0272_),
    .A2(_0276_),
    .A3(_0283_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1997_ (.I0(_1083_),
    .I1(_1096_),
    .S(_0951_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1998_ (.A1(_0286_),
    .A2(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1999_ (.A1(\mod.pc[4] ),
    .A2(_0281_),
    .B(_0267_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2000_ (.A1(_0281_),
    .A2(_0288_),
    .B(_0289_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2001_ (.A1(_0272_),
    .A2(_0276_),
    .A3(_0283_),
    .A4(_0287_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2002_ (.A1(\mod.pc[5] ),
    .A2(_1017_),
    .B(_1127_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2003_ (.A1(_0290_),
    .A2(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2004_ (.A1(_0290_),
    .A2(_0291_),
    .B(_0263_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2005_ (.I(_0223_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2006_ (.A1(_1118_),
    .A2(_0262_),
    .B1(_0292_),
    .B2(_0293_),
    .C(_0294_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2007_ (.I(_0241_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2008_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2009_ (.I(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2010_ (.I(_0241_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2011_ (.I(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2012_ (.A1(\mod.pc_1[0] ),
    .A2(_0299_),
    .B(_0267_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2013_ (.A1(_0781_),
    .A2(_0297_),
    .B(_0300_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2014_ (.I(_0266_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2015_ (.A1(\mod.pc_1[1] ),
    .A2(_0299_),
    .B(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2016_ (.A1(_0269_),
    .A2(_0297_),
    .B(_0302_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2017_ (.A1(\mod.pc_1[2] ),
    .A2(_0299_),
    .B(_0301_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2018_ (.A1(_1013_),
    .A2(_0297_),
    .B(_0303_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2019_ (.A1(\mod.pc_1[3] ),
    .A2(_0299_),
    .B(_0301_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2020_ (.A1(_0282_),
    .A2(_0297_),
    .B(_0304_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2021_ (.I(_0296_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2022_ (.I(_0298_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2023_ (.A1(\mod.pc_1[4] ),
    .A2(_0306_),
    .B(_0301_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2024_ (.A1(_1083_),
    .A2(_0305_),
    .B(_0307_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2025_ (.I(_0221_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2026_ (.I(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2027_ (.A1(\mod.pc_1[5] ),
    .A2(_0306_),
    .B(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2028_ (.A1(_1118_),
    .A2(_0305_),
    .B(_0310_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2029_ (.I(\mod.instr[0] ),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2030_ (.I(_0242_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2031_ (.I(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2032_ (.A1(\mod.des.des_dout[0] ),
    .A2(_0243_),
    .B(_0309_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2033_ (.A1(_0311_),
    .A2(_0313_),
    .B(_0314_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2034_ (.I(\mod.instr[1] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2035_ (.A1(\mod.des.des_dout[1] ),
    .A2(_0243_),
    .B(_0309_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2036_ (.A1(_0315_),
    .A2(_0313_),
    .B(_0316_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2037_ (.I(\mod.instr[2] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2038_ (.A1(\mod.des.des_dout[2] ),
    .A2(_0243_),
    .B(_0309_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2039_ (.A1(_0317_),
    .A2(_0313_),
    .B(_0318_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2040_ (.I(\mod.instr[3] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2041_ (.I(_0242_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2042_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2043_ (.I(_0308_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2044_ (.A1(\mod.des.des_dout[3] ),
    .A2(_0321_),
    .B(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2045_ (.A1(_0319_),
    .A2(_0313_),
    .B(_0323_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2046_ (.I(\mod.instr[4] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2047_ (.I(_0312_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2048_ (.A1(\mod.des.des_dout[4] ),
    .A2(_0321_),
    .B(_0322_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2049_ (.A1(_0324_),
    .A2(_0325_),
    .B(_0326_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2050_ (.I(\mod.instr[5] ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2051_ (.A1(\mod.des.des_dout[5] ),
    .A2(_0321_),
    .B(_0322_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2052_ (.A1(_0327_),
    .A2(_0325_),
    .B(_0328_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2053_ (.I(\mod.instr[6] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2054_ (.A1(\mod.des.des_dout[6] ),
    .A2(_0321_),
    .B(_0322_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2055_ (.A1(_0329_),
    .A2(_0325_),
    .B(_0330_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2056_ (.I(\mod.instr[7] ),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2057_ (.I(_0320_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2058_ (.I(_0308_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2059_ (.A1(\mod.des.des_dout[7] ),
    .A2(_0332_),
    .B(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2060_ (.A1(_0331_),
    .A2(_0325_),
    .B(_0334_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2061_ (.I(\mod.instr[8] ),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2062_ (.I(_0312_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2063_ (.A1(\mod.des.des_dout[8] ),
    .A2(_0332_),
    .B(_0333_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2064_ (.A1(_0335_),
    .A2(_0336_),
    .B(_0337_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2065_ (.I(\mod.instr[9] ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2066_ (.A1(\mod.des.des_dout[9] ),
    .A2(_0332_),
    .B(_0333_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2067_ (.A1(_0338_),
    .A2(_0336_),
    .B(_0339_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2068_ (.I(\mod.instr[10] ),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2069_ (.A1(\mod.des.des_dout[10] ),
    .A2(_0332_),
    .B(_0333_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2070_ (.A1(_0340_),
    .A2(_0336_),
    .B(_0341_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2071_ (.I(\mod.instr[11] ),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2072_ (.I(_0320_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2073_ (.I(_0308_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2074_ (.A1(\mod.des.des_dout[11] ),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2075_ (.A1(_0342_),
    .A2(_0336_),
    .B(_0345_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2076_ (.I(\mod.instr[12] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2077_ (.I(_0320_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2078_ (.A1(\mod.des.des_dout[12] ),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2079_ (.A1(_0346_),
    .A2(_0347_),
    .B(_0348_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2080_ (.I(\mod.instr[13] ),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2081_ (.A1(\mod.des.des_dout[13] ),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2082_ (.A1(_0349_),
    .A2(_0347_),
    .B(_0350_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2083_ (.I(\mod.instr[14] ),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2084_ (.A1(\mod.des.des_dout[14] ),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2085_ (.A1(_0351_),
    .A2(_0347_),
    .B(_0352_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2086_ (.I(\mod.instr[15] ),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2087_ (.A1(\mod.des.des_dout[15] ),
    .A2(_0312_),
    .B(_0222_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2088_ (.A1(_0353_),
    .A2(_0347_),
    .B(_0354_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2089_ (.A1(\mod.valid1 ),
    .A2(_0241_),
    .A3(_0229_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2090_ (.I(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2091_ (.A1(_0539_),
    .A2(_0228_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2092_ (.A1(_0356_),
    .A2(_0357_),
    .B(_0246_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2093_ (.I(_0295_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2094_ (.I(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2095_ (.A1(_0631_),
    .A2(_0359_),
    .B1(_0356_),
    .B2(\mod.instr[0] ),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2096_ (.A1(_0225_),
    .A2(_0360_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2097_ (.I(_0224_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2098_ (.A1(_0800_),
    .A2(_0359_),
    .B1(_0356_),
    .B2(\mod.instr[1] ),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2099_ (.A1(_0361_),
    .A2(_0362_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2100_ (.A1(_0776_),
    .A2(_0359_),
    .B1(_0356_),
    .B2(\mod.instr[2] ),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2101_ (.A1(_0361_),
    .A2(_0363_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2102_ (.I(_0355_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2103_ (.I(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2104_ (.A1(_0806_),
    .A2(_0359_),
    .B1(_0365_),
    .B2(\mod.instr[3] ),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2105_ (.A1(_0361_),
    .A2(_0366_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2106_ (.I(_0808_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2107_ (.I(_0358_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2108_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0365_),
    .B2(\mod.instr[4] ),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2109_ (.A1(_0361_),
    .A2(_0369_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2110_ (.I(_0224_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2111_ (.I(\mod.instr_2[5] ),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2112_ (.A1(_0371_),
    .A2(_0368_),
    .B1(_0365_),
    .B2(\mod.instr[5] ),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2113_ (.A1(_0370_),
    .A2(_0372_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2114_ (.A1(_0996_),
    .A2(_0368_),
    .B1(_0365_),
    .B2(\mod.instr[6] ),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2115_ (.A1(_0370_),
    .A2(_0373_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2116_ (.I(_0364_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2117_ (.A1(_1072_),
    .A2(_0368_),
    .B1(_0374_),
    .B2(\mod.instr[7] ),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2118_ (.A1(_0370_),
    .A2(_0375_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2119_ (.I(_0358_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2120_ (.A1(_0769_),
    .A2(_0376_),
    .B1(_0374_),
    .B2(\mod.instr[8] ),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2121_ (.A1(_0370_),
    .A2(_0377_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2122_ (.I(_0224_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2123_ (.A1(_0783_),
    .A2(_0376_),
    .B1(_0374_),
    .B2(\mod.instr[9] ),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2124_ (.A1(_0378_),
    .A2(_0379_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2125_ (.A1(_0787_),
    .A2(_0376_),
    .B1(_0374_),
    .B2(\mod.instr[10] ),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2126_ (.A1(_0378_),
    .A2(_0380_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2127_ (.I(_0364_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2128_ (.A1(_0577_),
    .A2(_0376_),
    .B1(_0381_),
    .B2(\mod.instr[11] ),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2129_ (.A1(_0378_),
    .A2(_0382_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2130_ (.I(_0298_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2131_ (.A1(_0696_),
    .A2(_0383_),
    .B1(_0381_),
    .B2(\mod.instr[12] ),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2132_ (.A1(_0378_),
    .A2(_0384_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2133_ (.A1(_0693_),
    .A2(_0383_),
    .B1(_0381_),
    .B2(\mod.instr[13] ),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2134_ (.A1(_0232_),
    .A2(_0385_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2135_ (.A1(\mod.instr_2[14] ),
    .A2(_0383_),
    .B1(_0381_),
    .B2(\mod.instr[14] ),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2136_ (.A1(_0232_),
    .A2(_0386_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2137_ (.A1(_0545_),
    .A2(_0383_),
    .B1(_0364_),
    .B2(\mod.instr[15] ),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2138_ (.A1(_0232_),
    .A2(_0387_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2139_ (.I(_0227_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2140_ (.A1(\mod.pc_1[0] ),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2141_ (.I(_0295_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2142_ (.A1(\mod.pc_2[0] ),
    .A2(_0390_),
    .B(_0003_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2143_ (.A1(_0389_),
    .A2(_0391_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2144_ (.A1(\mod.pc_1[1] ),
    .A2(_0388_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2145_ (.A1(_0953_),
    .A2(_0390_),
    .B(_0003_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2146_ (.A1(_0392_),
    .A2(_0393_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2147_ (.A1(\mod.pc_1[2] ),
    .A2(_0388_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2148_ (.A1(_1019_),
    .A2(_0390_),
    .B(_0003_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2149_ (.A1(_0394_),
    .A2(_0395_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2150_ (.A1(\mod.pc_1[3] ),
    .A2(_0388_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2151_ (.I(_0358_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2152_ (.I(_0266_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2153_ (.A1(_1051_),
    .A2(_0397_),
    .B(_0398_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2154_ (.A1(_0396_),
    .A2(_0399_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2155_ (.A1(\mod.pc_1[4] ),
    .A2(_0244_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2156_ (.A1(\mod.pc_2[4] ),
    .A2(_0397_),
    .B(_0398_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2157_ (.A1(_0400_),
    .A2(_0401_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2158_ (.A1(\mod.pc_1[5] ),
    .A2(_0244_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2159_ (.A1(\mod.pc_2[5] ),
    .A2(_0397_),
    .B(_0398_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2160_ (.A1(_0402_),
    .A2(_0403_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2161_ (.A1(_0539_),
    .A2(_0295_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2162_ (.A1(_0247_),
    .A2(\mod.ins_ldr_3 ),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2163_ (.A1(\mod.valid_out3 ),
    .A2(_0244_),
    .A3(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2164_ (.A1(_0404_),
    .A2(_0406_),
    .B(_0246_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2165_ (.I(_0804_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2166_ (.A1(_0407_),
    .A2(_0885_),
    .B(_0404_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2167_ (.A1(_0939_),
    .A2(_0404_),
    .B(_0408_),
    .C(_0280_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2168_ (.A1(\mod.ri_3 ),
    .A2(_0296_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2169_ (.A1(_0713_),
    .A2(_0390_),
    .B(_0409_),
    .C(_0280_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2170_ (.A1(_0407_),
    .A2(_0298_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2171_ (.A1(\mod.ins_ldr_3 ),
    .A2(_0228_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2172_ (.A1(_0410_),
    .A2(_0411_),
    .B(_0246_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2173_ (.A1(\mod.rd_3[0] ),
    .A2(_0306_),
    .B(_0222_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2174_ (.A1(_0813_),
    .A2(_0305_),
    .B(_0412_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(\mod.rd_3[1] ),
    .A2(_0397_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2176_ (.A1(_0367_),
    .A2(_0228_),
    .B(_0398_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2177_ (.A1(_0413_),
    .A2(_0414_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2178_ (.A1(\mod.rd_3[2] ),
    .A2(_0306_),
    .B(_0222_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2179_ (.A1(_1159_),
    .A2(_0305_),
    .B(_0415_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2180_ (.A1(_0249_),
    .A2(_0223_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2181_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2182_ (.A1(_0782_),
    .A2(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2183_ (.I(_0418_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2184_ (.A1(_0407_),
    .A2(_0810_),
    .A3(_0296_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(\mod.ldr_hzd[1] ),
    .A2(_0417_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2186_ (.A1(_0371_),
    .A2(_0252_),
    .A3(_0419_),
    .B(_0420_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2187_ (.A1(_0367_),
    .A2(_0407_),
    .A3(_1014_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(_0813_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2189_ (.A1(_0247_),
    .A2(_1159_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2190_ (.I(_0416_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2191_ (.A1(_0795_),
    .A2(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2192_ (.A1(_0280_),
    .A2(_0422_),
    .A3(_0423_),
    .B(_0425_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(_0806_),
    .A2(_0421_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2194_ (.A1(\mod.ldr_hzd[3] ),
    .A2(_0424_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2195_ (.A1(_0294_),
    .A2(_0423_),
    .A3(_0426_),
    .B(_0427_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2196_ (.A1(_0371_),
    .A2(_0266_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2197_ (.A1(_0367_),
    .A2(_0806_),
    .A3(_0410_),
    .A4(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2198_ (.A1(\mod.ldr_hzd[4] ),
    .A2(_0417_),
    .B(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2199_ (.I(_0430_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2200_ (.A1(\mod.ldr_hzd[5] ),
    .A2(_0417_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2201_ (.A1(_0419_),
    .A2(_0428_),
    .B(_0431_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2202_ (.A1(_0247_),
    .A2(_0371_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_0424_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2204_ (.A1(_0294_),
    .A2(_0422_),
    .A3(_0432_),
    .B(_0433_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(\mod.ldr_hzd[7] ),
    .A2(_0424_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2206_ (.A1(_0294_),
    .A2(_0426_),
    .A3(_0432_),
    .B(_0434_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2207_ (.A1(\mod.des.des_counter[2] ),
    .A2(_0532_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2208_ (.I(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2209_ (.I0(\mod.des.des_dout[12] ),
    .I1(net1),
    .S(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2210_ (.I(_0437_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2211_ (.I0(\mod.des.des_dout[13] ),
    .I1(net2),
    .S(_0436_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2212_ (.I(_0438_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2213_ (.I0(\mod.des.des_dout[14] ),
    .I1(net3),
    .S(_0435_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2214_ (.I(_0439_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2215_ (.I0(\mod.des.des_dout[15] ),
    .I1(net4),
    .S(_0435_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_0440_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2217_ (.A1(net5),
    .A2(_0436_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2218_ (.A1(_0188_),
    .A2(_0436_),
    .B(_0441_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2219_ (.I0(\mod.des.des_dout[17] ),
    .I1(net6),
    .S(_0435_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2220_ (.I(_0442_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2221_ (.A1(_1152_),
    .A2(_1156_),
    .A3(_1164_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2222_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2223_ (.I0(_0192_),
    .I1(\mod.registers.r7[0] ),
    .S(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2224_ (.I(_0445_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2225_ (.I(_0443_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2226_ (.I(_0443_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2227_ (.A1(\mod.registers.r7[1] ),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2228_ (.A1(_0202_),
    .A2(_0446_),
    .B(_0448_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2229_ (.A1(\mod.registers.r7[2] ),
    .A2(_0447_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2230_ (.A1(_0209_),
    .A2(_0446_),
    .B(_0449_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2231_ (.I0(_0215_),
    .I1(\mod.registers.r7[3] ),
    .S(_0444_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2232_ (.I(_0450_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(\mod.registers.r7[4] ),
    .A2(_0447_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2234_ (.A1(_0165_),
    .A2(_0446_),
    .B(_0451_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2235_ (.I0(_0173_),
    .I1(\mod.registers.r7[5] ),
    .S(_0444_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2236_ (.I(_0452_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2237_ (.A1(\mod.registers.r7[6] ),
    .A2(_0447_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2238_ (.A1(_0182_),
    .A2(_0446_),
    .B(_0453_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2239_ (.I0(_0186_),
    .I1(\mod.registers.r7[7] ),
    .S(_0444_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2240_ (.I(_0454_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2241_ (.A1(_0534_),
    .A2(_1029_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2242_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2243_ (.I0(\mod.des.des_dout[0] ),
    .I1(net1),
    .S(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2244_ (.I(_0457_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2245_ (.I0(\mod.des.des_dout[1] ),
    .I1(net2),
    .S(_0456_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2246_ (.I(_0458_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2247_ (.I0(\mod.des.des_dout[2] ),
    .I1(net3),
    .S(_0456_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2248_ (.I(_0459_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2249_ (.I0(\mod.des.des_dout[3] ),
    .I1(net4),
    .S(_0456_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2250_ (.I(_0460_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2251_ (.I0(\mod.des.des_dout[4] ),
    .I1(net5),
    .S(_0455_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2252_ (.I(_0461_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2253_ (.I0(\mod.des.des_dout[5] ),
    .I1(net6),
    .S(_0455_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2254_ (.I(_0462_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2255_ (.A1(_0534_),
    .A2(_0531_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2256_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2257_ (.I0(\mod.des.des_dout[6] ),
    .I1(net1),
    .S(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2258_ (.I(_0465_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2259_ (.I0(\mod.des.des_dout[7] ),
    .I1(net2),
    .S(_0464_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2260_ (.I(_0466_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2261_ (.I0(\mod.des.des_dout[8] ),
    .I1(net3),
    .S(_0464_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2262_ (.I(_0467_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2263_ (.I0(\mod.des.des_dout[9] ),
    .I1(net4),
    .S(_0464_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2264_ (.I(_0468_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2265_ (.I0(\mod.des.des_dout[10] ),
    .I1(net5),
    .S(_0463_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2266_ (.I(_0469_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2267_ (.I0(\mod.des.des_dout[11] ),
    .I1(net6),
    .S(_0463_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2268_ (.I(_0470_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2269_ (.I(_0225_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2270_ (.A1(_1159_),
    .A2(_1154_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2271_ (.A1(\mod.rd_3[2] ),
    .A2(_1154_),
    .B(_0471_),
    .C(_1163_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2272_ (.A1(_1158_),
    .A2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2273_ (.I(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2274_ (.I(_0473_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2275_ (.A1(_0191_),
    .A2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2276_ (.A1(_0695_),
    .A2(_0474_),
    .B(_0476_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2277_ (.I(_0473_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2278_ (.A1(\mod.registers.r1[1] ),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2279_ (.A1(_0202_),
    .A2(_0474_),
    .B(_0478_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2280_ (.A1(\mod.registers.r1[2] ),
    .A2(_0477_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2281_ (.A1(_0209_),
    .A2(_0474_),
    .B(_0479_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2282_ (.I0(_0215_),
    .I1(\mod.registers.r1[3] ),
    .S(_0475_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2283_ (.I(_0480_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2284_ (.A1(\mod.registers.r1[4] ),
    .A2(_0477_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2285_ (.A1(_0165_),
    .A2(_0474_),
    .B(_0481_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2286_ (.I0(_0173_),
    .I1(\mod.registers.r1[5] ),
    .S(_0475_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2287_ (.I(_0482_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2288_ (.A1(\mod.registers.r1[6] ),
    .A2(_0475_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2289_ (.A1(_0182_),
    .A2(_0477_),
    .B(_0483_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2290_ (.I0(_0186_),
    .I1(\mod.registers.r1[7] ),
    .S(_0473_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2291_ (.I(_0484_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2292_ (.A1(_0194_),
    .A2(_0472_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2293_ (.I(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2294_ (.I0(_0192_),
    .I1(\mod.registers.r2[0] ),
    .S(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2295_ (.I(_0487_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2296_ (.I(_0485_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2297_ (.I(_0485_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2298_ (.A1(\mod.registers.r2[1] ),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2299_ (.A1(_0201_),
    .A2(_0488_),
    .B(_0490_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(\mod.registers.r2[2] ),
    .A2(_0489_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2301_ (.A1(_0208_),
    .A2(_0488_),
    .B(_0491_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2302_ (.I0(_0215_),
    .I1(\mod.registers.r2[3] ),
    .S(_0486_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2303_ (.I(_0492_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2304_ (.A1(\mod.registers.r2[4] ),
    .A2(_0489_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2305_ (.A1(_0164_),
    .A2(_0488_),
    .B(_0493_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2306_ (.I0(_0172_),
    .I1(\mod.registers.r2[5] ),
    .S(_0486_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2307_ (.I(_0494_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2308_ (.A1(\mod.registers.r2[6] ),
    .A2(_0489_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2309_ (.A1(_0181_),
    .A2(_0488_),
    .B(_0495_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2310_ (.I0(_0185_),
    .I1(\mod.registers.r2[7] ),
    .S(_0486_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2311_ (.I(_0496_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2312_ (.A1(_1152_),
    .A2(_1156_),
    .A3(_0472_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2313_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2314_ (.I0(_0192_),
    .I1(\mod.registers.r3[0] ),
    .S(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2315_ (.I(_0499_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2316_ (.I(_0497_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2317_ (.I(_0497_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2318_ (.A1(\mod.registers.r3[1] ),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2319_ (.A1(_0201_),
    .A2(_0500_),
    .B(_0502_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2320_ (.A1(\mod.registers.r3[2] ),
    .A2(_0501_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2321_ (.A1(_0208_),
    .A2(_0500_),
    .B(_0503_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2322_ (.I0(_0214_),
    .I1(\mod.registers.r3[3] ),
    .S(_0498_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2323_ (.I(_0504_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(\mod.registers.r3[4] ),
    .A2(_0501_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2325_ (.A1(_0164_),
    .A2(_0500_),
    .B(_0505_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2326_ (.I0(_0172_),
    .I1(\mod.registers.r3[5] ),
    .S(_0498_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2327_ (.I(_0506_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2328_ (.A1(\mod.registers.r3[6] ),
    .A2(_0501_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2329_ (.A1(_0181_),
    .A2(_0500_),
    .B(_0507_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2330_ (.I0(_0185_),
    .I1(\mod.registers.r3[7] ),
    .S(_0498_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2331_ (.I(_0508_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2332_ (.A1(_0193_),
    .A2(_1157_),
    .A3(_1164_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2333_ (.I(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2334_ (.I0(_0191_),
    .I1(\mod.registers.r4[0] ),
    .S(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2335_ (.I(_0511_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2336_ (.I(_0509_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2337_ (.I(_0509_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2338_ (.A1(\mod.registers.r4[1] ),
    .A2(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2339_ (.A1(_0201_),
    .A2(_0512_),
    .B(_0514_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2340_ (.A1(\mod.registers.r4[2] ),
    .A2(_0513_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2341_ (.A1(_0208_),
    .A2(_0512_),
    .B(_0515_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2342_ (.I0(_0214_),
    .I1(\mod.registers.r4[3] ),
    .S(_0510_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2343_ (.I(_0516_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2344_ (.A1(\mod.registers.r4[4] ),
    .A2(_0513_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2345_ (.A1(_0164_),
    .A2(_0512_),
    .B(_0517_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2346_ (.I0(_0172_),
    .I1(\mod.registers.r4[5] ),
    .S(_0510_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2347_ (.I(_0518_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2348_ (.A1(\mod.registers.r4[6] ),
    .A2(_0513_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2349_ (.A1(_0181_),
    .A2(_0512_),
    .B(_0519_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2350_ (.I0(_0185_),
    .I1(\mod.registers.r4[7] ),
    .S(_0510_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2351_ (.I(_0520_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2352_ (.I0(_0191_),
    .I1(\mod.registers.r5[0] ),
    .S(_0174_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2353_ (.I(_0521_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2354_ (.A1(\mod.registers.r5[1] ),
    .A2(_0166_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2355_ (.A1(_1166_),
    .A2(_0202_),
    .B(_0522_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2356_ (.A1(\mod.registers.r5[2] ),
    .A2(_0166_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2357_ (.A1(_1166_),
    .A2(_0209_),
    .B(_0523_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2358_ (.I0(_0214_),
    .I1(\mod.registers.r5[3] ),
    .S(_0174_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2359_ (.I(_0524_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2360_ (.D(_0007_),
    .CLK(net60),
    .Q(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2361_ (.D(_0008_),
    .CLK(net73),
    .Q(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2362_ (.D(_0009_),
    .CLK(net59),
    .Q(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2363_ (.D(_0010_),
    .CLK(net73),
    .Q(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2364_ (.D(_0011_),
    .CLK(net70),
    .Q(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2365_ (.D(_0012_),
    .CLK(net55),
    .Q(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2366_ (.D(_0013_),
    .CLK(net55),
    .Q(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2367_ (.D(_0014_),
    .CLK(net59),
    .Q(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2368_ (.D(_0015_),
    .CLK(net60),
    .Q(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2369_ (.D(_0016_),
    .CLK(net71),
    .Q(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2370_ (.D(_0017_),
    .CLK(net60),
    .Q(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2371_ (.D(_0018_),
    .CLK(net69),
    .Q(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2372_ (.D(_0000_),
    .SETN(_0003_),
    .CLK(net83),
    .Q(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2373_ (.D(_0001_),
    .SETN(_0004_),
    .CLK(net83),
    .Q(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2374_ (.D(_0002_),
    .SETN(_0005_),
    .CLK(net81),
    .Q(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2375_ (.D(_0019_),
    .CLK(net19),
    .Q(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2376_ (.D(_0020_),
    .CLK(net86),
    .Q(\mod.des.des_dout[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2377_ (.D(_0021_),
    .CLK(net84),
    .Q(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2378_ (.D(_0022_),
    .CLK(net85),
    .Q(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2379_ (.D(_0023_),
    .CLK(net86),
    .Q(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2380_ (.D(_0024_),
    .CLK(net84),
    .Q(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2381_ (.D(_0025_),
    .CLK(net88),
    .Q(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2382_ (.D(_0026_),
    .CLK(net19),
    .Q(\mod.valid1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2383_ (.D(_0027_),
    .CLK(net43),
    .Q(\mod.pc0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2384_ (.D(_0028_),
    .CLK(net41),
    .Q(\mod.pc0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2385_ (.D(_0029_),
    .CLK(net43),
    .Q(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2386_ (.D(_0030_),
    .CLK(net40),
    .Q(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2387_ (.D(_0031_),
    .CLK(net40),
    .Q(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2388_ (.D(_0032_),
    .CLK(net40),
    .Q(\mod.pc0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2389_ (.D(_0033_),
    .CLK(net39),
    .Q(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2390_ (.D(_0034_),
    .CLK(net41),
    .Q(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2391_ (.D(_0035_),
    .CLK(net39),
    .Q(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2392_ (.D(_0036_),
    .CLK(net39),
    .Q(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2393_ (.D(_0037_),
    .CLK(net39),
    .Q(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2394_ (.D(_0038_),
    .CLK(net40),
    .Q(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2395_ (.D(_0039_),
    .CLK(net35),
    .Q(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2396_ (.D(_0040_),
    .CLK(net35),
    .Q(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2397_ (.D(_0041_),
    .CLK(net34),
    .Q(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2398_ (.D(_0042_),
    .CLK(net34),
    .Q(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2399_ (.D(_0043_),
    .CLK(net33),
    .Q(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2400_ (.D(_0044_),
    .CLK(net34),
    .Q(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2401_ (.D(_0045_),
    .CLK(net19),
    .Q(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2402_ (.D(_0046_),
    .CLK(net18),
    .Q(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2403_ (.D(_0047_),
    .CLK(net18),
    .Q(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2404_ (.D(_0048_),
    .CLK(net18),
    .Q(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2405_ (.D(_0049_),
    .CLK(net18),
    .Q(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2406_ (.D(_0050_),
    .CLK(net26),
    .Q(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2407_ (.D(_0051_),
    .CLK(net26),
    .Q(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2408_ (.D(_0052_),
    .CLK(net26),
    .Q(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2409_ (.D(_0053_),
    .CLK(net27),
    .Q(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2410_ (.D(_0054_),
    .CLK(net27),
    .Q(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2411_ (.D(_0055_),
    .CLK(net27),
    .Q(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2412_ (.D(_0056_),
    .CLK(net27),
    .Q(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2413_ (.D(_0057_),
    .CLK(net45),
    .Q(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2414_ (.D(_0058_),
    .CLK(net45),
    .Q(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2415_ (.D(_0059_),
    .CLK(net45),
    .Q(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2416_ (.D(_0060_),
    .CLK(net28),
    .Q(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2417_ (.D(_0061_),
    .CLK(net36),
    .Q(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2418_ (.D(_0062_),
    .CLK(net30),
    .Q(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2419_ (.D(_0063_),
    .CLK(net30),
    .Q(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2420_ (.D(_0064_),
    .CLK(net31),
    .Q(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2421_ (.D(_0065_),
    .CLK(net25),
    .Q(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2422_ (.D(_0066_),
    .CLK(net30),
    .Q(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2423_ (.D(_0067_),
    .CLK(net29),
    .Q(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2424_ (.D(_0068_),
    .CLK(net28),
    .Q(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2425_ (.D(_0069_),
    .CLK(net28),
    .Q(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2426_ (.D(_0070_),
    .CLK(net29),
    .Q(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2427_ (.D(_0071_),
    .CLK(net46),
    .Q(\mod.instr_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2428_ (.D(_0072_),
    .CLK(net46),
    .Q(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2429_ (.D(_0073_),
    .CLK(net45),
    .Q(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2430_ (.D(_0074_),
    .CLK(net50),
    .Q(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2431_ (.D(_0075_),
    .CLK(net50),
    .Q(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2432_ (.D(_0076_),
    .CLK(net50),
    .Q(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2433_ (.D(_0077_),
    .CLK(net50),
    .Q(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2434_ (.D(_0078_),
    .CLK(net37),
    .Q(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2435_ (.D(_0079_),
    .CLK(net36),
    .Q(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2436_ (.D(_0080_),
    .CLK(net37),
    .Q(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2437_ (.D(_0081_),
    .CLK(net33),
    .Q(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2438_ (.D(_0082_),
    .CLK(net33),
    .Q(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2439_ (.D(_0083_),
    .CLK(net33),
    .Q(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2440_ (.D(_0084_),
    .CLK(net23),
    .Q(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2441_ (.D(_0085_),
    .CLK(net36),
    .Q(\mod.des.des_din[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2442_ (.D(_0086_),
    .CLK(net36),
    .Q(\mod.ri_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2443_ (.D(_0087_),
    .CLK(net21),
    .Q(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2444_ (.D(_0088_),
    .CLK(net23),
    .Q(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2445_ (.D(_0089_),
    .CLK(net21),
    .Q(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2446_ (.D(_0090_),
    .CLK(net22),
    .Q(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2447_ (.D(_0091_),
    .CLK(net30),
    .Q(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2448_ (.D(_0092_),
    .CLK(net22),
    .Q(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2449_ (.D(_0093_),
    .CLK(net20),
    .Q(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2450_ (.D(_0094_),
    .CLK(net20),
    .Q(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2451_ (.D(_0095_),
    .CLK(net22),
    .Q(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2452_ (.D(_0096_),
    .CLK(net22),
    .Q(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2453_ (.D(_0097_),
    .CLK(net20),
    .Q(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2454_ (.D(_0098_),
    .CLK(net20),
    .Q(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2455_ (.D(_0099_),
    .CLK(net87),
    .Q(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2456_ (.D(_0100_),
    .CLK(net84),
    .Q(\mod.des.des_dout[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2457_ (.D(_0101_),
    .CLK(net85),
    .Q(\mod.des.des_dout[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2458_ (.D(_0102_),
    .CLK(net79),
    .Q(\mod.des.des_dout[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2459_ (.D(_0103_),
    .CLK(net84),
    .Q(\mod.des.des_dout[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2460_ (.D(_0104_),
    .CLK(net88),
    .Q(\mod.des.des_dout[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2461_ (.D(_0105_),
    .CLK(net70),
    .Q(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2462_ (.D(_0106_),
    .CLK(net54),
    .Q(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2463_ (.D(_0107_),
    .CLK(net54),
    .Q(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2464_ (.D(_0108_),
    .CLK(net58),
    .Q(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2465_ (.D(_0109_),
    .CLK(net60),
    .Q(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2466_ (.D(_0110_),
    .CLK(net69),
    .Q(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2467_ (.D(_0111_),
    .CLK(net58),
    .Q(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2468_ (.D(_0112_),
    .CLK(net69),
    .Q(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2469_ (.D(_0113_),
    .CLK(net77),
    .Q(\mod.des.des_dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2470_ (.D(_0114_),
    .CLK(net77),
    .Q(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2471_ (.D(_0115_),
    .CLK(net77),
    .Q(\mod.des.des_dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2472_ (.D(_0116_),
    .CLK(net77),
    .Q(\mod.des.des_dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2473_ (.D(_0117_),
    .CLK(net78),
    .Q(\mod.des.des_dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2474_ (.D(_0118_),
    .CLK(net79),
    .Q(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2475_ (.D(_0119_),
    .CLK(net79),
    .Q(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2476_ (.D(_0120_),
    .CLK(net79),
    .Q(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2477_ (.D(_0121_),
    .CLK(net80),
    .Q(\mod.des.des_dout[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2478_ (.D(_0122_),
    .CLK(net80),
    .Q(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2479_ (.D(_0123_),
    .CLK(net87),
    .Q(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2480_ (.D(_0124_),
    .CLK(net87),
    .Q(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2481_ (.D(_0125_),
    .RN(_0006_),
    .CLK(net81),
    .Q(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2482_ (.D(_0126_),
    .CLK(net72),
    .Q(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2483_ (.D(_0127_),
    .CLK(net53),
    .Q(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2484_ (.D(_0128_),
    .CLK(net53),
    .Q(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2485_ (.D(_0129_),
    .CLK(net58),
    .Q(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2486_ (.D(_0130_),
    .CLK(net62),
    .Q(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2487_ (.D(_0131_),
    .CLK(net69),
    .Q(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2488_ (.D(_0132_),
    .CLK(net62),
    .Q(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2489_ (.D(_0133_),
    .CLK(net72),
    .Q(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2490_ (.D(_0134_),
    .CLK(net65),
    .Q(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2491_ (.D(_0135_),
    .CLK(net47),
    .Q(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2492_ (.D(_0136_),
    .CLK(net51),
    .Q(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2493_ (.D(_0137_),
    .CLK(net58),
    .Q(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2494_ (.D(_0138_),
    .CLK(net51),
    .Q(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2495_ (.D(_0139_),
    .CLK(net68),
    .Q(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2496_ (.D(_0140_),
    .CLK(net51),
    .Q(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2497_ (.D(_0141_),
    .CLK(net66),
    .Q(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2498_ (.D(_0142_),
    .CLK(net65),
    .Q(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2499_ (.D(_0143_),
    .CLK(net48),
    .Q(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2500_ (.D(_0144_),
    .CLK(net47),
    .Q(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2501_ (.D(_0145_),
    .CLK(net65),
    .Q(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2502_ (.D(_0146_),
    .CLK(net47),
    .Q(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2503_ (.D(_0147_),
    .CLK(net66),
    .Q(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2504_ (.D(_0148_),
    .CLK(net47),
    .Q(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2505_ (.D(_0149_),
    .CLK(net66),
    .Q(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2506_ (.D(_0150_),
    .CLK(net65),
    .Q(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2507_ (.D(_0151_),
    .CLK(net48),
    .Q(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2508_ (.D(_0152_),
    .CLK(net57),
    .Q(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2509_ (.D(_0153_),
    .CLK(net51),
    .Q(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2510_ (.D(_0154_),
    .CLK(net53),
    .Q(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2511_ (.D(_0155_),
    .CLK(net74),
    .Q(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2512_ (.D(_0156_),
    .CLK(net53),
    .Q(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2513_ (.D(_0157_),
    .CLK(net73),
    .Q(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2514_ (.D(_0158_),
    .CLK(net70),
    .Q(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2515_ (.D(_0159_),
    .CLK(net54),
    .Q(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2516_ (.D(_0160_),
    .CLK(net54),
    .Q(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2517_ (.D(_0161_),
    .CLK(net70),
    .Q(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout18 (.I(net19),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout19 (.I(net25),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout20 (.I(net24),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout21 (.I(net24),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout22 (.I(net24),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout23 (.I(net24),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout24 (.I(net25),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout25 (.I(net32),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout26 (.I(net29),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout27 (.I(net28),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout28 (.I(net29),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout29 (.I(net31),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout32 (.I(net44),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(net38),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout35 (.I(net38),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout36 (.I(net38),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout38 (.I(net42),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net41),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net43),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net76),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net49),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net49),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net52),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net52),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net64),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net57),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net56),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net63),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net61),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout60 (.I(net62),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net63),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net75),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout65 (.I(net67),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net74),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout69 (.I(net71),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net72),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net74),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net76),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(\mod.clk ),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net82),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout79 (.I(net81),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net89),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net8),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__B2 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__SETN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__SETN (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__RN (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__D (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__D (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__D (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__D (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__B2 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__I (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A1 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__B (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__I0 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__I0 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I0 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A3 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__I (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A2 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__I0 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__I0 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__I0 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__I (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__B (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__B1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I0 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__I0 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A1 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__I (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I0 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__I0 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I0 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__I0 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A2 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__S (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__S (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__S (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__S (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__B (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__I (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__B (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__I0 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__I0 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__I0 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__B (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__B (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__B (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__I (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__I (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__I (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__I (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__I (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__I (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__I (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__I (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__I (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A2 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__B (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__S (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__S (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__I (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__S (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__S (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__S (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__S (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A2 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__I (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__I (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__I (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__I (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__B (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__B (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__B (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__B (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__I (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__I (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__I (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__C (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__C (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__C (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__C (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__C (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__C (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__C (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__B (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__C (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__C (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__C (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__C (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I0 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__C (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A3 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__I (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__B (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__B (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__B (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__B (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__B (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__B (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__B (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__B (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__B (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__B1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__B1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__B1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__B (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A4 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__B (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__S (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__S (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__S (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__S (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__S (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__S (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__S (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__S (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__S (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__S (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__S (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__S (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__S (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__S (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__S (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A3 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__S (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__S (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__S (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__S (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__S (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__S (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__S (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__B (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__B (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__S (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__S (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__S (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__S (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1181__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1194__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__B (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1297__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1286__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1336__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__S (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1258__I (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__I (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1332__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1316__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__B1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__B1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__B1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__B1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__B1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1318__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__C1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__C1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__I (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__B1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__C1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__C1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__C1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1224__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1227__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1227__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__A3 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__A3 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A3 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1227__A3 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__C (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__B (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__B1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__B1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__B1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1236__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__B1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__C1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__B1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1240__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__B1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__B1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__B1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1290__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__A3 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A3 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__A3 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__B1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__C1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__C1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__I (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__C2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__B1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__C2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__B1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__C2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__B1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__B1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__B1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__B1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__B1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__B1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1251__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__B1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__B (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1337__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1261__I (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1391__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1278__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1270__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__B1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__C1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1365__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1276__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__B2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1304__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1288__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1288__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A3 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A3 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1303__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__S0 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__I1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A3 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__A3 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1294__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1330__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__S (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1302__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__I (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1313__B (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__I0 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__I1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__I (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A3 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A3 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__C (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1353__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1353__A3 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__B2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__B (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__C (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__B2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A3 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A3 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A3 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__C (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1427__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__I (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__B (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__C (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1429__I (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__B (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__B (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__B (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__B2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__I (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__B (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__I1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__C (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__C (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__C (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__B (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__A3 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__B2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A3 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__C (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__B (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1503__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__B (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1539__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__B (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__C (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__I (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__B1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__B1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__B2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__A2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__B (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__I1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__B (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A3 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__C (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__B (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__B (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__B2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__S (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__B1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__B (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__S (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A3 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__B (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__B (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A3 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A3 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A3 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__B2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__I0 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A3 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__B1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__B2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__B2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__B2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__B (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__B2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__C (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__I0 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__B1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__I0 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__B (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__B1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__I1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__B1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__B (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__B (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__B (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A3 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A3 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__C (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__B1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__B1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A4 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__B (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__B (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__S (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__I (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__B (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__I (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__S (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__B (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__B (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__C (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__C (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A3 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A3 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A3 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__B1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__I (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__I (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__A1 (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__I0 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__I0 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__I0 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__I0 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__A1 (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1330__A1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__B (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1292__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A2 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B2 (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__B2 (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__I (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__B2 (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__I (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__B2 (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__I (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__B2 (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__I (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__B2 (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__I (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__B2 (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__I (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__B2 (.I(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__I (.I(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__B2 (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__I (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__B2 (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__I (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__B2 (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__I (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A1 (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A1 (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1215__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__I1 (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__I0 (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1300__I1 (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__A1 (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1200__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1310__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A1 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A3 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A1 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1439__I (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__I (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A1 (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A1 (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A1 (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__B2 (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__I (.I(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A1 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A4 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__B2 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I0 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A3 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__A1 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I1 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A2 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I2 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A1 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A1 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A1 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I3 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__I (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__I1 (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__I (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__I (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__I0 (.I(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A1 (.I(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__I (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1319__A3 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__B2 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__I1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__I1 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__B2 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__B2 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__I1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__B2 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__I1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__A3 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__C1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1332__A3 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1317__A3 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__B2 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__I1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__B2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I1 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A3 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__A1 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A3 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__B2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1318__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__I1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__C2 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__A1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__C2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__C2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__I1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__A1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__C2 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__B2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__C2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__I1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__B2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__C2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__B2 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__B2 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__B2 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__I1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__B2 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__I1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__B2 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__C1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__C2 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__I1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__C2 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__B2 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__I1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__C1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__B2 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__I1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__I1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__I1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__CLK (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__CLK (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1043 ();
 assign io_oeb[0] = net90;
 assign io_oeb[10] = net100;
 assign io_oeb[11] = net101;
 assign io_oeb[12] = net102;
 assign io_oeb[13] = net103;
 assign io_oeb[14] = net104;
 assign io_oeb[15] = net105;
 assign io_oeb[16] = net106;
 assign io_oeb[17] = net107;
 assign io_oeb[18] = net108;
 assign io_oeb[19] = net109;
 assign io_oeb[1] = net91;
 assign io_oeb[20] = net110;
 assign io_oeb[21] = net111;
 assign io_oeb[22] = net112;
 assign io_oeb[23] = net113;
 assign io_oeb[24] = net114;
 assign io_oeb[25] = net115;
 assign io_oeb[26] = net116;
 assign io_oeb[27] = net117;
 assign io_oeb[28] = net118;
 assign io_oeb[29] = net119;
 assign io_oeb[2] = net92;
 assign io_oeb[30] = net120;
 assign io_oeb[31] = net121;
 assign io_oeb[32] = net122;
 assign io_oeb[33] = net123;
 assign io_oeb[34] = net124;
 assign io_oeb[35] = net125;
 assign io_oeb[36] = net126;
 assign io_oeb[37] = net127;
 assign io_oeb[3] = net93;
 assign io_oeb[4] = net94;
 assign io_oeb[5] = net95;
 assign io_oeb[6] = net96;
 assign io_oeb[7] = net97;
 assign io_oeb[8] = net98;
 assign io_oeb[9] = net99;
 assign io_out[0] = net128;
 assign io_out[10] = net138;
 assign io_out[11] = net139;
 assign io_out[12] = net140;
 assign io_out[13] = net141;
 assign io_out[14] = net142;
 assign io_out[15] = net143;
 assign io_out[16] = net144;
 assign io_out[1] = net129;
 assign io_out[25] = net145;
 assign io_out[26] = net146;
 assign io_out[27] = net147;
 assign io_out[28] = net148;
 assign io_out[29] = net149;
 assign io_out[2] = net130;
 assign io_out[30] = net150;
 assign io_out[31] = net151;
 assign io_out[32] = net152;
 assign io_out[33] = net153;
 assign io_out[34] = net154;
 assign io_out[35] = net155;
 assign io_out[36] = net156;
 assign io_out[37] = net157;
 assign io_out[3] = net131;
 assign io_out[4] = net132;
 assign io_out[5] = net133;
 assign io_out[6] = net134;
 assign io_out[7] = net135;
 assign io_out[8] = net136;
 assign io_out[9] = net137;
 assign la_data_out[0] = net158;
 assign la_data_out[10] = net168;
 assign la_data_out[11] = net169;
 assign la_data_out[12] = net170;
 assign la_data_out[13] = net171;
 assign la_data_out[14] = net172;
 assign la_data_out[15] = net173;
 assign la_data_out[16] = net174;
 assign la_data_out[17] = net175;
 assign la_data_out[18] = net176;
 assign la_data_out[19] = net177;
 assign la_data_out[1] = net159;
 assign la_data_out[20] = net178;
 assign la_data_out[21] = net179;
 assign la_data_out[22] = net180;
 assign la_data_out[23] = net181;
 assign la_data_out[24] = net182;
 assign la_data_out[25] = net183;
 assign la_data_out[26] = net184;
 assign la_data_out[27] = net185;
 assign la_data_out[28] = net186;
 assign la_data_out[29] = net187;
 assign la_data_out[2] = net160;
 assign la_data_out[30] = net188;
 assign la_data_out[31] = net189;
 assign la_data_out[32] = net190;
 assign la_data_out[33] = net191;
 assign la_data_out[34] = net192;
 assign la_data_out[35] = net193;
 assign la_data_out[36] = net194;
 assign la_data_out[37] = net195;
 assign la_data_out[38] = net196;
 assign la_data_out[39] = net197;
 assign la_data_out[3] = net161;
 assign la_data_out[40] = net198;
 assign la_data_out[41] = net199;
 assign la_data_out[42] = net200;
 assign la_data_out[43] = net201;
 assign la_data_out[44] = net202;
 assign la_data_out[45] = net203;
 assign la_data_out[46] = net204;
 assign la_data_out[47] = net205;
 assign la_data_out[48] = net206;
 assign la_data_out[49] = net207;
 assign la_data_out[4] = net162;
 assign la_data_out[50] = net208;
 assign la_data_out[51] = net209;
 assign la_data_out[52] = net210;
 assign la_data_out[53] = net211;
 assign la_data_out[54] = net212;
 assign la_data_out[55] = net213;
 assign la_data_out[56] = net214;
 assign la_data_out[57] = net215;
 assign la_data_out[58] = net216;
 assign la_data_out[59] = net217;
 assign la_data_out[5] = net163;
 assign la_data_out[60] = net218;
 assign la_data_out[61] = net219;
 assign la_data_out[62] = net220;
 assign la_data_out[63] = net221;
 assign la_data_out[6] = net164;
 assign la_data_out[7] = net165;
 assign la_data_out[8] = net166;
 assign la_data_out[9] = net167;
 assign user_irq[0] = net222;
 assign user_irq[1] = net223;
 assign user_irq[2] = net224;
 assign wbs_ack_o = net225;
 assign wbs_dat_o[0] = net226;
 assign wbs_dat_o[10] = net236;
 assign wbs_dat_o[11] = net237;
 assign wbs_dat_o[12] = net238;
 assign wbs_dat_o[13] = net239;
 assign wbs_dat_o[14] = net240;
 assign wbs_dat_o[15] = net241;
 assign wbs_dat_o[16] = net242;
 assign wbs_dat_o[17] = net243;
 assign wbs_dat_o[18] = net244;
 assign wbs_dat_o[19] = net245;
 assign wbs_dat_o[1] = net227;
 assign wbs_dat_o[20] = net246;
 assign wbs_dat_o[21] = net247;
 assign wbs_dat_o[22] = net248;
 assign wbs_dat_o[23] = net249;
 assign wbs_dat_o[24] = net250;
 assign wbs_dat_o[25] = net251;
 assign wbs_dat_o[26] = net252;
 assign wbs_dat_o[27] = net253;
 assign wbs_dat_o[28] = net254;
 assign wbs_dat_o[29] = net255;
 assign wbs_dat_o[2] = net228;
 assign wbs_dat_o[30] = net256;
 assign wbs_dat_o[31] = net257;
 assign wbs_dat_o[3] = net229;
 assign wbs_dat_o[4] = net230;
 assign wbs_dat_o[5] = net231;
 assign wbs_dat_o[6] = net232;
 assign wbs_dat_o[7] = net233;
 assign wbs_dat_o[8] = net234;
 assign wbs_dat_o[9] = net235;
endmodule

