// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire net152;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net153;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net154;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net191;
 wire net192;
 wire net190;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net212;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net213;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net214;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net215;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net216;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire \mod.clk ;
 wire \mod.des.des_counter[0] ;
 wire \mod.des.des_counter[1] ;
 wire \mod.des.des_counter[2] ;
 wire \mod.des.des_dout[0] ;
 wire \mod.des.des_dout[10] ;
 wire \mod.des.des_dout[11] ;
 wire \mod.des.des_dout[12] ;
 wire \mod.des.des_dout[13] ;
 wire \mod.des.des_dout[14] ;
 wire \mod.des.des_dout[15] ;
 wire \mod.des.des_dout[16] ;
 wire \mod.des.des_dout[17] ;
 wire \mod.des.des_dout[18] ;
 wire \mod.des.des_dout[19] ;
 wire \mod.des.des_dout[1] ;
 wire \mod.des.des_dout[20] ;
 wire \mod.des.des_dout[21] ;
 wire \mod.des.des_dout[22] ;
 wire \mod.des.des_dout[23] ;
 wire \mod.des.des_dout[24] ;
 wire \mod.des.des_dout[25] ;
 wire \mod.des.des_dout[26] ;
 wire \mod.des.des_dout[27] ;
 wire \mod.des.des_dout[28] ;
 wire \mod.des.des_dout[29] ;
 wire \mod.des.des_dout[2] ;
 wire \mod.des.des_dout[30] ;
 wire \mod.des.des_dout[31] ;
 wire \mod.des.des_dout[32] ;
 wire \mod.des.des_dout[33] ;
 wire \mod.des.des_dout[3] ;
 wire \mod.des.des_dout[4] ;
 wire \mod.des.des_dout[5] ;
 wire \mod.des.des_dout[6] ;
 wire \mod.des.des_dout[7] ;
 wire \mod.des.des_dout[8] ;
 wire \mod.des.des_dout[9] ;
 wire \mod.funct3[0] ;
 wire \mod.funct3[1] ;
 wire \mod.funct3[2] ;
 wire \mod.funct7[0] ;
 wire \mod.funct7[1] ;
 wire \mod.funct7[2] ;
 wire \mod.ins_ldr_3 ;
 wire \mod.instr[0] ;
 wire \mod.instr[10] ;
 wire \mod.instr[11] ;
 wire \mod.instr[12] ;
 wire \mod.instr[13] ;
 wire \mod.instr[14] ;
 wire \mod.instr[15] ;
 wire \mod.instr[16] ;
 wire \mod.instr[17] ;
 wire \mod.instr[1] ;
 wire \mod.instr[2] ;
 wire \mod.instr[3] ;
 wire \mod.instr[4] ;
 wire \mod.instr[5] ;
 wire \mod.instr[6] ;
 wire \mod.instr[7] ;
 wire \mod.instr[8] ;
 wire \mod.instr[9] ;
 wire \mod.instr_2[0] ;
 wire \mod.instr_2[10] ;
 wire \mod.instr_2[11] ;
 wire \mod.instr_2[12] ;
 wire \mod.instr_2[13] ;
 wire \mod.instr_2[14] ;
 wire \mod.instr_2[1] ;
 wire \mod.instr_2[2] ;
 wire \mod.instr_2[3] ;
 wire \mod.instr_2[4] ;
 wire \mod.instr_2[5] ;
 wire \mod.instr_2[9] ;
 wire \mod.ldr_hzd[0] ;
 wire \mod.ldr_hzd[1] ;
 wire \mod.ldr_hzd[2] ;
 wire \mod.ldr_hzd[3] ;
 wire \mod.ldr_hzd[4] ;
 wire \mod.ldr_hzd[5] ;
 wire \mod.ldr_hzd[6] ;
 wire \mod.ldr_hzd[7] ;
 wire \mod.pc0[0] ;
 wire \mod.pc0[10] ;
 wire \mod.pc0[11] ;
 wire \mod.pc0[12] ;
 wire \mod.pc0[13] ;
 wire \mod.pc0[1] ;
 wire \mod.pc0[2] ;
 wire \mod.pc0[3] ;
 wire \mod.pc0[4] ;
 wire \mod.pc0[5] ;
 wire \mod.pc0[6] ;
 wire \mod.pc0[7] ;
 wire \mod.pc0[8] ;
 wire \mod.pc0[9] ;
 wire \mod.pc[0] ;
 wire \mod.pc[10] ;
 wire \mod.pc[11] ;
 wire \mod.pc[12] ;
 wire \mod.pc[13] ;
 wire \mod.pc[1] ;
 wire \mod.pc[2] ;
 wire \mod.pc[3] ;
 wire \mod.pc[4] ;
 wire \mod.pc[5] ;
 wire \mod.pc[6] ;
 wire \mod.pc[7] ;
 wire \mod.pc[8] ;
 wire \mod.pc[9] ;
 wire \mod.pc_1[0] ;
 wire \mod.pc_1[10] ;
 wire \mod.pc_1[11] ;
 wire \mod.pc_1[12] ;
 wire \mod.pc_1[13] ;
 wire \mod.pc_1[1] ;
 wire \mod.pc_1[2] ;
 wire \mod.pc_1[3] ;
 wire \mod.pc_1[4] ;
 wire \mod.pc_1[5] ;
 wire \mod.pc_1[6] ;
 wire \mod.pc_1[7] ;
 wire \mod.pc_1[8] ;
 wire \mod.pc_1[9] ;
 wire \mod.pc_2[0] ;
 wire \mod.pc_2[10] ;
 wire \mod.pc_2[11] ;
 wire \mod.pc_2[12] ;
 wire \mod.pc_2[13] ;
 wire \mod.pc_2[1] ;
 wire \mod.pc_2[2] ;
 wire \mod.pc_2[3] ;
 wire \mod.pc_2[4] ;
 wire \mod.pc_2[5] ;
 wire \mod.pc_2[6] ;
 wire \mod.pc_2[7] ;
 wire \mod.pc_2[8] ;
 wire \mod.pc_2[9] ;
 wire \mod.rd_3[0] ;
 wire \mod.rd_3[1] ;
 wire \mod.rd_3[2] ;
 wire \mod.registers.r1[0] ;
 wire \mod.registers.r1[10] ;
 wire \mod.registers.r1[11] ;
 wire \mod.registers.r1[12] ;
 wire \mod.registers.r1[13] ;
 wire \mod.registers.r1[14] ;
 wire \mod.registers.r1[15] ;
 wire \mod.registers.r1[1] ;
 wire \mod.registers.r1[2] ;
 wire \mod.registers.r1[3] ;
 wire \mod.registers.r1[4] ;
 wire \mod.registers.r1[5] ;
 wire \mod.registers.r1[6] ;
 wire \mod.registers.r1[7] ;
 wire \mod.registers.r1[8] ;
 wire \mod.registers.r1[9] ;
 wire \mod.registers.r2[0] ;
 wire \mod.registers.r2[10] ;
 wire \mod.registers.r2[11] ;
 wire \mod.registers.r2[12] ;
 wire \mod.registers.r2[13] ;
 wire \mod.registers.r2[14] ;
 wire \mod.registers.r2[15] ;
 wire \mod.registers.r2[1] ;
 wire \mod.registers.r2[2] ;
 wire \mod.registers.r2[3] ;
 wire \mod.registers.r2[4] ;
 wire \mod.registers.r2[5] ;
 wire \mod.registers.r2[6] ;
 wire \mod.registers.r2[7] ;
 wire \mod.registers.r2[8] ;
 wire \mod.registers.r2[9] ;
 wire \mod.registers.r3[0] ;
 wire \mod.registers.r3[10] ;
 wire \mod.registers.r3[11] ;
 wire \mod.registers.r3[12] ;
 wire \mod.registers.r3[13] ;
 wire \mod.registers.r3[14] ;
 wire \mod.registers.r3[15] ;
 wire \mod.registers.r3[1] ;
 wire \mod.registers.r3[2] ;
 wire \mod.registers.r3[3] ;
 wire \mod.registers.r3[4] ;
 wire \mod.registers.r3[5] ;
 wire \mod.registers.r3[6] ;
 wire \mod.registers.r3[7] ;
 wire \mod.registers.r3[8] ;
 wire \mod.registers.r3[9] ;
 wire \mod.registers.r4[0] ;
 wire \mod.registers.r4[10] ;
 wire \mod.registers.r4[11] ;
 wire \mod.registers.r4[12] ;
 wire \mod.registers.r4[13] ;
 wire \mod.registers.r4[14] ;
 wire \mod.registers.r4[15] ;
 wire \mod.registers.r4[1] ;
 wire \mod.registers.r4[2] ;
 wire \mod.registers.r4[3] ;
 wire \mod.registers.r4[4] ;
 wire \mod.registers.r4[5] ;
 wire \mod.registers.r4[6] ;
 wire \mod.registers.r4[7] ;
 wire \mod.registers.r4[8] ;
 wire \mod.registers.r4[9] ;
 wire \mod.registers.r5[0] ;
 wire \mod.registers.r5[10] ;
 wire \mod.registers.r5[11] ;
 wire \mod.registers.r5[12] ;
 wire \mod.registers.r5[13] ;
 wire \mod.registers.r5[14] ;
 wire \mod.registers.r5[15] ;
 wire \mod.registers.r5[1] ;
 wire \mod.registers.r5[2] ;
 wire \mod.registers.r5[3] ;
 wire \mod.registers.r5[4] ;
 wire \mod.registers.r5[5] ;
 wire \mod.registers.r5[6] ;
 wire \mod.registers.r5[7] ;
 wire \mod.registers.r5[8] ;
 wire \mod.registers.r5[9] ;
 wire \mod.registers.r6[0] ;
 wire \mod.registers.r6[10] ;
 wire \mod.registers.r6[11] ;
 wire \mod.registers.r6[12] ;
 wire \mod.registers.r6[13] ;
 wire \mod.registers.r6[14] ;
 wire \mod.registers.r6[15] ;
 wire \mod.registers.r6[1] ;
 wire \mod.registers.r6[2] ;
 wire \mod.registers.r6[3] ;
 wire \mod.registers.r6[4] ;
 wire \mod.registers.r6[5] ;
 wire \mod.registers.r6[6] ;
 wire \mod.registers.r6[7] ;
 wire \mod.registers.r6[8] ;
 wire \mod.registers.r6[9] ;
 wire \mod.registers.r7[0] ;
 wire \mod.registers.r7[10] ;
 wire \mod.registers.r7[11] ;
 wire \mod.registers.r7[12] ;
 wire \mod.registers.r7[13] ;
 wire \mod.registers.r7[14] ;
 wire \mod.registers.r7[15] ;
 wire \mod.registers.r7[1] ;
 wire \mod.registers.r7[2] ;
 wire \mod.registers.r7[3] ;
 wire \mod.registers.r7[4] ;
 wire \mod.registers.r7[5] ;
 wire \mod.registers.r7[6] ;
 wire \mod.registers.r7[7] ;
 wire \mod.registers.r7[8] ;
 wire \mod.registers.r7[9] ;
 wire \mod.ri_3 ;
 wire \mod.valid0 ;
 wire \mod.valid1 ;
 wire \mod.valid2 ;
 wire \mod.valid_out3 ;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net280;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net281;
 wire net309;
 wire net310;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2551_ (.I(\mod.instr[10] ),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2552_ (.A1(\mod.des.des_dout[10] ),
    .A2(_1962_),
    .B(_1963_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2553_ (.A1(_1965_),
    .A2(_1959_),
    .B(_1966_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2554_ (.I(\mod.instr[11] ),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2555_ (.A1(\mod.des.des_dout[11] ),
    .A2(_1962_),
    .B(_1963_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2556_ (.A1(_1967_),
    .A2(_1959_),
    .B(_1968_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2557_ (.I(\mod.instr[12] ),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2558_ (.I(_1924_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2559_ (.A1(\mod.des.des_dout[12] ),
    .A2(_1962_),
    .B(_1963_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2560_ (.A1(_1969_),
    .A2(_1970_),
    .B(_1971_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2561_ (.I(\mod.instr[13] ),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2562_ (.I(_1923_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2563_ (.I(_1508_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2564_ (.A1(\mod.des.des_dout[13] ),
    .A2(_1973_),
    .B(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2565_ (.A1(_1972_),
    .A2(_1970_),
    .B(_1975_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2566_ (.I(\mod.instr[14] ),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2567_ (.A1(\mod.des.des_dout[14] ),
    .A2(_1973_),
    .B(_1974_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2568_ (.A1(_1976_),
    .A2(_1970_),
    .B(_1977_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2569_ (.I(\mod.instr[15] ),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2570_ (.A1(\mod.des.des_dout[15] ),
    .A2(_1973_),
    .B(_1974_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2571_ (.A1(_1978_),
    .A2(_1970_),
    .B(_1979_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2572_ (.I(\mod.instr[16] ),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2573_ (.A1(\mod.des.des_dout[16] ),
    .A2(_1973_),
    .B(_1974_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2574_ (.A1(_1980_),
    .A2(_1925_),
    .B(_1981_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2575_ (.I(\mod.instr[17] ),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2576_ (.A1(\mod.des.des_dout[17] ),
    .A2(_1936_),
    .B(_1509_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2577_ (.A1(_1982_),
    .A2(_1925_),
    .B(_1983_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2578_ (.A1(_0003_),
    .A2(_1315_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2579_ (.I(_1984_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2580_ (.A1(_1854_),
    .A2(_1354_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2581_ (.A1(_1854_),
    .A2(_1368_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2582_ (.I(_1853_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2583_ (.A1(_1985_),
    .A2(_1395_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2584_ (.A1(_1985_),
    .A2(_1422_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2585_ (.A1(_1985_),
    .A2(_1458_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2586_ (.A1(_0003_),
    .A2(_1481_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2587_ (.I(_1986_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2588_ (.A1(_1985_),
    .A2(_1295_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2589_ (.I(_1853_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2590_ (.A1(_1987_),
    .A2(_1337_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2591_ (.A1(_1987_),
    .A2(_1383_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2592_ (.A1(_1987_),
    .A2(_1409_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2593_ (.A1(_1425_),
    .A2(_1433_),
    .B(_1815_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2594_ (.A1(_1987_),
    .A2(_1449_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2595_ (.I(_1793_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2596_ (.I(_1988_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2597_ (.A1(_1989_),
    .A2(_1474_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2598_ (.I(_1812_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2599_ (.A1(\mod.pc_1[0] ),
    .A2(_1990_),
    .B1(_1933_),
    .B2(\mod.pc_2[0] ),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2600_ (.I(_1991_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2601_ (.A1(\mod.pc_1[1] ),
    .A2(_1990_),
    .B1(_1933_),
    .B2(\mod.pc_2[1] ),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2602_ (.I(_1992_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2603_ (.A1(\mod.pc_1[2] ),
    .A2(_1990_),
    .B1(_1933_),
    .B2(_1264_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2604_ (.I(_1993_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2605_ (.I(_1931_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2606_ (.A1(\mod.pc_1[3] ),
    .A2(_1990_),
    .B1(_1994_),
    .B2(\mod.pc_2[3] ),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2607_ (.I(_1995_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2608_ (.I(_1812_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2609_ (.A1(\mod.pc_1[4] ),
    .A2(_1996_),
    .B1(_1994_),
    .B2(_1260_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2610_ (.I(_1997_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2611_ (.A1(\mod.pc_1[5] ),
    .A2(_1996_),
    .B1(_1994_),
    .B2(_1257_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2612_ (.I(_1998_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2613_ (.A1(\mod.pc_1[6] ),
    .A2(_1996_),
    .B1(_1994_),
    .B2(_1254_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2614_ (.I(_1999_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2615_ (.I(_1931_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2616_ (.A1(\mod.pc_1[7] ),
    .A2(_1996_),
    .B1(_2000_),
    .B2(_1252_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2617_ (.I(_2001_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2618_ (.I(_1812_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2619_ (.A1(\mod.pc_1[8] ),
    .A2(_2002_),
    .B1(_2000_),
    .B2(_1327_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2620_ (.I(_2003_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2621_ (.A1(\mod.pc_1[9] ),
    .A2(_2002_),
    .B1(_2000_),
    .B2(_1373_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2622_ (.I(_2004_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2623_ (.A1(\mod.pc_1[10] ),
    .A2(_2002_),
    .B1(_2000_),
    .B2(_1399_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2624_ (.I(_2005_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2625_ (.A1(\mod.pc_1[11] ),
    .A2(_2002_),
    .B1(_1932_),
    .B2(_1438_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2626_ (.I(_2006_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2627_ (.A1(\mod.pc_1[12] ),
    .A2(_1813_),
    .B1(_1932_),
    .B2(_1464_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2628_ (.I(_2007_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2629_ (.A1(\mod.pc_1[13] ),
    .A2(_1813_),
    .B1(_1932_),
    .B2(\mod.pc_2[13] ),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2630_ (.I(_2008_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2631_ (.A1(_2128_),
    .A2(_1797_),
    .B1(_1930_),
    .B2(\mod.instr[0] ),
    .C(_1809_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2632_ (.I(_2009_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2633_ (.I(_1929_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2634_ (.I(_2010_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2635_ (.A1(_1204_),
    .A2(_1808_),
    .B1(_2011_),
    .B2(\mod.instr[1] ),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2636_ (.A1(_1989_),
    .A2(_2012_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2637_ (.A1(_2125_),
    .A2(_1797_),
    .B1(_1930_),
    .B2(\mod.instr[2] ),
    .C(_1809_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2638_ (.I(_2013_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2639_ (.A1(_1227_),
    .A2(_1808_),
    .B1(_2011_),
    .B2(\mod.instr[3] ),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2640_ (.A1(_1989_),
    .A2(_2014_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2641_ (.I(_1796_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2642_ (.A1(_1230_),
    .A2(_2015_),
    .B1(_2011_),
    .B2(\mod.instr[4] ),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2643_ (.A1(_1989_),
    .A2(_2016_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2644_ (.I(_1988_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2645_ (.A1(_1510_),
    .A2(_2015_),
    .B1(_2011_),
    .B2(\mod.instr[5] ),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2646_ (.A1(_2017_),
    .A2(_2018_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2647_ (.I(_1929_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2648_ (.A1(_0738_),
    .A2(_2015_),
    .B1(_2019_),
    .B2(\mod.instr[6] ),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_2017_),
    .A2(_2020_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2650_ (.A1(_0645_),
    .A2(_2015_),
    .B1(_2019_),
    .B2(\mod.instr[7] ),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2651_ (.A1(_2017_),
    .A2(_2021_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2652_ (.A1(_0820_),
    .A2(_1797_),
    .B1(_1930_),
    .B2(\mod.instr[8] ),
    .C(_1809_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2653_ (.I(_2022_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2654_ (.I(_1796_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2655_ (.A1(_2164_),
    .A2(_2023_),
    .B1(_2019_),
    .B2(\mod.instr[9] ),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2656_ (.A1(_2017_),
    .A2(_2024_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2657_ (.I(_1988_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2658_ (.A1(_2154_),
    .A2(_2023_),
    .B1(_2019_),
    .B2(\mod.instr[10] ),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2659_ (.A1(_2025_),
    .A2(_2026_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2660_ (.I(_1929_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2661_ (.A1(_2181_),
    .A2(_2023_),
    .B1(_2027_),
    .B2(\mod.instr[11] ),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2662_ (.A1(_2025_),
    .A2(_2028_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2663_ (.A1(_1216_),
    .A2(_2023_),
    .B1(_2027_),
    .B2(\mod.instr[12] ),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2664_ (.A1(_2025_),
    .A2(_2029_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2665_ (.I(_1424_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2666_ (.A1(_0428_),
    .A2(_2030_),
    .B1(_2027_),
    .B2(\mod.instr[13] ),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2667_ (.A1(_2025_),
    .A2(_2031_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2668_ (.I(_1988_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2669_ (.A1(_0423_),
    .A2(_2030_),
    .B1(_2027_),
    .B2(\mod.instr[14] ),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2670_ (.A1(_2032_),
    .A2(_2033_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2671_ (.A1(\mod.funct7[0] ),
    .A2(_2030_),
    .B1(_2010_),
    .B2(\mod.instr[15] ),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2672_ (.A1(_2032_),
    .A2(_2034_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2673_ (.A1(_2243_),
    .A2(_2030_),
    .B1(_2010_),
    .B2(\mod.instr[16] ),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2674_ (.A1(_2032_),
    .A2(_2035_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2675_ (.A1(_1437_),
    .A2(_1823_),
    .B1(_2010_),
    .B2(\mod.instr[17] ),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2676_ (.A1(_2032_),
    .A2(_2036_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2677_ (.A1(\mod.valid2 ),
    .A2(_1823_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2678_ (.A1(\mod.valid_out3 ),
    .A2(_1814_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2679_ (.A1(_2037_),
    .A2(_2038_),
    .B(_1815_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2680_ (.A1(_1510_),
    .A2(_1224_),
    .A3(_1813_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2681_ (.A1(_1234_),
    .A2(_2039_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2682_ (.A1(_1226_),
    .A2(_1227_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2683_ (.A1(_1224_),
    .A2(_1807_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2684_ (.A1(_2040_),
    .A2(_2041_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(_1230_),
    .A2(_1232_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2686_ (.A1(_2042_),
    .A2(_2041_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2687_ (.A1(_1234_),
    .A2(_2041_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2688_ (.A1(_1230_),
    .A2(_1227_),
    .A3(_2039_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2689_ (.A1(_2040_),
    .A2(_2039_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2690_ (.A1(_2042_),
    .A2(_2039_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2691_ (.A1(\mod.des.des_counter[2] ),
    .A2(\mod.des.des_counter[1] ),
    .A3(\mod.des.des_counter[0] ),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2692_ (.I(_2043_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2693_ (.I0(\mod.des.des_dout[0] ),
    .I1(net13),
    .S(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2694_ (.I(_2045_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2695_ (.I0(\mod.des.des_dout[1] ),
    .I1(net14),
    .S(_2044_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2696_ (.I(_2046_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2697_ (.I0(\mod.des.des_dout[2] ),
    .I1(net15),
    .S(_2044_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2698_ (.I(_2047_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2699_ (.I0(\mod.des.des_dout[3] ),
    .I1(net16),
    .S(_2044_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_2048_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2701_ (.I(_2043_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2702_ (.I0(\mod.des.des_dout[4] ),
    .I1(net17),
    .S(_2049_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2703_ (.I(_2050_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2704_ (.I0(\mod.des.des_dout[5] ),
    .I1(net18),
    .S(_2049_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2705_ (.I(_2051_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2706_ (.I0(\mod.des.des_dout[6] ),
    .I1(net2),
    .S(_2049_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2707_ (.I(_2052_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2708_ (.I0(\mod.des.des_dout[7] ),
    .I1(net3),
    .S(_2049_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2709_ (.I(_2053_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2710_ (.I(_2043_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2711_ (.I0(\mod.des.des_dout[8] ),
    .I1(net4),
    .S(_2054_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2712_ (.I(_2055_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2713_ (.I0(\mod.des.des_dout[9] ),
    .I1(net5),
    .S(_2054_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2714_ (.I(_2056_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2715_ (.I0(\mod.des.des_dout[10] ),
    .I1(net6),
    .S(_2054_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2716_ (.I(_2057_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2717_ (.I0(\mod.des.des_dout[11] ),
    .I1(net7),
    .S(_2054_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2718_ (.I(_2058_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2719_ (.I(_2043_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2720_ (.I0(\mod.des.des_dout[12] ),
    .I1(net8),
    .S(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2721_ (.I(_2060_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2722_ (.I0(\mod.des.des_dout[13] ),
    .I1(net9),
    .S(_2059_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2723_ (.I(_2061_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2724_ (.I0(\mod.des.des_dout[14] ),
    .I1(net10),
    .S(_2059_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2725_ (.I(_2062_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2726_ (.I0(\mod.des.des_dout[15] ),
    .I1(net11),
    .S(_2059_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2727_ (.I(_2063_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2728_ (.A1(_1517_),
    .A2(_1522_),
    .A3(_1715_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2729_ (.I(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2730_ (.I(_2065_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2731_ (.I0(_1660_),
    .I1(\mod.registers.r7[0] ),
    .S(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2732_ (.I(_2067_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_2065_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2734_ (.I(_2064_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(\mod.registers.r7[1] ),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2736_ (.A1(_1550_),
    .A2(_2068_),
    .B(_2070_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2737_ (.A1(\mod.registers.r7[2] ),
    .A2(_2069_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2738_ (.A1(_1559_),
    .A2(_2068_),
    .B(_2071_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2739_ (.A1(\mod.registers.r7[3] ),
    .A2(_2069_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2740_ (.A1(_1565_),
    .A2(_2068_),
    .B(_2072_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2741_ (.A1(\mod.registers.r7[4] ),
    .A2(_2069_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2742_ (.A1(_1570_),
    .A2(_2068_),
    .B(_2073_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2743_ (.I0(_1580_),
    .I1(\mod.registers.r7[5] ),
    .S(_2066_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2744_ (.I(_2074_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2745_ (.I0(_1594_),
    .I1(\mod.registers.r7[6] ),
    .S(_2066_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2746_ (.I(_2075_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2747_ (.I0(_1601_),
    .I1(\mod.registers.r7[7] ),
    .S(_2066_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2748_ (.I(_2076_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2749_ (.I(_2065_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2750_ (.I0(_1610_),
    .I1(\mod.registers.r7[8] ),
    .S(_2077_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2751_ (.I(_2078_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2752_ (.I0(_1616_),
    .I1(\mod.registers.r7[9] ),
    .S(_2077_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2753_ (.I(_2079_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2754_ (.I0(_1624_),
    .I1(\mod.registers.r7[10] ),
    .S(_2077_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2755_ (.I(_2080_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2756_ (.I(_2065_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2757_ (.I(_2064_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2758_ (.A1(\mod.registers.r7[11] ),
    .A2(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2759_ (.A1(_1631_),
    .A2(_2081_),
    .B(_2083_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(\mod.registers.r7[12] ),
    .A2(_2082_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2761_ (.A1(_1638_),
    .A2(_2081_),
    .B(_2084_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2762_ (.A1(\mod.registers.r7[13] ),
    .A2(_2082_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2763_ (.A1(_1645_),
    .A2(_2081_),
    .B(_2085_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2764_ (.I0(_1652_),
    .I1(\mod.registers.r7[14] ),
    .S(_2077_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2765_ (.I(_2086_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2766_ (.A1(\mod.registers.r7[15] ),
    .A2(_2082_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2767_ (.A1(_1657_),
    .A2(_2081_),
    .B(_2087_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2768_ (.A1(\mod.des.des_counter[2] ),
    .A2(_1411_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2769_ (.I(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2770_ (.I(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2771_ (.I0(net13),
    .I1(\mod.des.des_dout[16] ),
    .S(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2772_ (.I(_2091_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2773_ (.I0(net14),
    .I1(\mod.des.des_dout[17] ),
    .S(_2090_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2774_ (.I(_2092_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2775_ (.A1(net15),
    .A2(_2090_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2776_ (.A1(_1539_),
    .A2(_2090_),
    .B(_2093_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2777_ (.I(_2089_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2778_ (.I0(net16),
    .I1(\mod.des.des_dout[19] ),
    .S(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2779_ (.I(_2095_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2780_ (.I0(net17),
    .I1(\mod.des.des_dout[20] ),
    .S(_2094_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2781_ (.I(_2096_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2782_ (.I0(net18),
    .I1(\mod.des.des_dout[21] ),
    .S(_2094_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2783_ (.I(_2097_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2784_ (.I0(net2),
    .I1(\mod.des.des_dout[22] ),
    .S(_2094_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2785_ (.I(_2098_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2786_ (.I(_2089_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2787_ (.I0(net3),
    .I1(\mod.des.des_dout[23] ),
    .S(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2788_ (.I(_2100_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2789_ (.I0(net4),
    .I1(\mod.des.des_dout[24] ),
    .S(_2099_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2790_ (.I(_2101_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2791_ (.I0(net5),
    .I1(\mod.des.des_dout[25] ),
    .S(_2099_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2792_ (.I(_2102_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2793_ (.I0(net6),
    .I1(\mod.des.des_dout[26] ),
    .S(_2099_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2794_ (.I(_2103_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2795_ (.I(_2088_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2796_ (.I0(net7),
    .I1(\mod.des.des_dout[27] ),
    .S(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2797_ (.I(_2105_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2798_ (.I0(net8),
    .I1(\mod.des.des_dout[28] ),
    .S(_2104_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2799_ (.I(_2106_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2800_ (.I0(net9),
    .I1(\mod.des.des_dout[29] ),
    .S(_2104_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2801_ (.I(_2107_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2802_ (.I0(net10),
    .I1(\mod.des.des_dout[30] ),
    .S(_2104_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2803_ (.I(_2108_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2804_ (.I0(net11),
    .I1(\mod.des.des_dout[31] ),
    .S(_2089_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2805_ (.I(_2109_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2806_ (.A1(\mod.des.des_counter[2] ),
    .A2(_2122_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2807_ (.A1(net13),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2808_ (.A1(_1648_),
    .A2(_2110_),
    .B(_2111_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2809_ (.I0(\mod.des.des_dout[33] ),
    .I1(net14),
    .S(_2110_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2810_ (.I(_2112_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2811_ (.I(\mod.des.des_counter[1] ),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2812_ (.I(\mod.des.des_counter[0] ),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2813_ (.A1(_2113_),
    .A2(_0000_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2814_ (.A1(net112),
    .A2(_2114_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2815_ (.I(_2115_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(_2113_),
    .A2(\mod.des.des_counter[0] ),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2817_ (.A1(\mod.des.des_counter[1] ),
    .A2(_0000_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2818_ (.A1(_2116_),
    .A2(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2819_ (.I(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2820_ (.I(_2119_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2821_ (.I(_2120_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2822_ (.A1(\mod.des.des_counter[2] ),
    .A2(_2114_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2823_ (.I(_2121_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2824_ (.A1(\mod.des.des_counter[1] ),
    .A2(_0000_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2825_ (.I(_2122_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2826_ (.I(\mod.instr_2[2] ),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2827_ (.I(_2124_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2828_ (.I(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2829_ (.I(\mod.instr_2[0] ),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2830_ (.I(_2127_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2831_ (.A1(_2126_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2832_ (.I(_2129_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2833_ (.I(\mod.instr_2[1] ),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2834_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_2131_),
    .A2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2836_ (.I(_2133_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2837_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2838_ (.I(_2135_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2839_ (.I(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2840_ (.I(\mod.instr_2[11] ),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2841_ (.I(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2842_ (.I(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2843_ (.I(_2140_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2844_ (.I(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2845_ (.I(\mod.instr_2[9] ),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2846_ (.A1(\mod.instr_2[10] ),
    .A2(_2143_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2847_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2848_ (.I(_2145_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2849_ (.A1(_2142_),
    .A2(_2146_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2850_ (.I(_2139_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2851_ (.I(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2852_ (.I(_2149_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2853_ (.I(\mod.instr_2[10] ),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2854_ (.I(_2151_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2855_ (.I(_2152_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2856_ (.I(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2857_ (.I(_2143_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2858_ (.I(_2155_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2859_ (.I(_2156_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2860_ (.A1(_2150_),
    .A2(_2154_),
    .A3(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2861_ (.A1(\mod.registers.r3[15] ),
    .A2(_2147_),
    .B1(_2158_),
    .B2(\mod.registers.r4[15] ),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2862_ (.I(\mod.instr_2[10] ),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2863_ (.I(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2864_ (.I(_2161_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2865_ (.I(_2162_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2866_ (.I(_2157_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2867_ (.A1(_2150_),
    .A2(_2163_),
    .A3(_2164_),
    .A4(\mod.registers.r1[15] ),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2868_ (.I(\mod.instr_2[11] ),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2869_ (.A1(_2166_),
    .A2(_2151_),
    .A3(_2143_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2870_ (.I(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2871_ (.I(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2872_ (.A1(\mod.registers.r7[15] ),
    .A2(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2873_ (.I(_2152_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2874_ (.I(_2171_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2875_ (.I(\mod.instr_2[9] ),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2876_ (.I(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2877_ (.I(_2174_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2878_ (.I(_2175_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2879_ (.I(_2176_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2880_ (.A1(_2150_),
    .A2(_2172_),
    .A3(_2177_),
    .A4(\mod.registers.r2[15] ),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2881_ (.I(_2166_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2882_ (.I(_2179_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2883_ (.I(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2884_ (.A1(_2181_),
    .A2(_2172_),
    .A3(_2177_),
    .A4(\mod.registers.r6[15] ),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2885_ (.A1(_2181_),
    .A2(_2163_),
    .A3(_2157_),
    .A4(\mod.registers.r5[15] ),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2886_ (.A1(_2178_),
    .A2(_2182_),
    .A3(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2887_ (.A1(_2159_),
    .A2(_2165_),
    .A3(_2170_),
    .A4(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2888_ (.A1(_2137_),
    .A2(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2889_ (.I(_2131_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2890_ (.A1(_2124_),
    .A2(_2127_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2891_ (.A1(_2187_),
    .A2(_2188_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2892_ (.I(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2893_ (.I(\mod.instr_2[14] ),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2894_ (.I(_2191_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2895_ (.I(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2896_ (.I(\mod.instr_2[13] ),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2897_ (.I(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2898_ (.I(_2195_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2899_ (.I(\mod.instr_2[12] ),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2900_ (.I(_2197_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2901_ (.I(_2198_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2902_ (.A1(_2193_),
    .A2(_2196_),
    .A3(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2903_ (.I(_2200_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2904_ (.I(\mod.instr_2[14] ),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2905_ (.I(_2202_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2906_ (.I(\mod.instr_2[13] ),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2907_ (.I(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2908_ (.I(\mod.instr_2[12] ),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2909_ (.I(_2206_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2910_ (.I(_2207_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2911_ (.A1(_2203_),
    .A2(_2205_),
    .A3(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2912_ (.I(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2913_ (.I(_2192_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2914_ (.I(_2204_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2915_ (.I(_2212_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2916_ (.I(_2207_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2917_ (.A1(_2211_),
    .A2(_2213_),
    .A3(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2918_ (.I(_2215_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2919_ (.A1(\mod.registers.r5[15] ),
    .A2(_2201_),
    .B1(_2210_),
    .B2(\mod.registers.r2[15] ),
    .C1(_2216_),
    .C2(\mod.registers.r6[15] ),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2920_ (.A1(_2202_),
    .A2(_2194_),
    .A3(_2206_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2921_ (.I(_2218_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2922_ (.I(_2219_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2923_ (.I(_2192_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2924_ (.A1(_2194_),
    .A2(_2206_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2925_ (.I(_2222_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2926_ (.A1(_2221_),
    .A2(_2223_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2927_ (.I(_2224_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2928_ (.A1(\mod.registers.r7[15] ),
    .A2(_2220_),
    .B1(_2225_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2929_ (.I(_2195_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2930_ (.A1(_2221_),
    .A2(_2227_),
    .A3(_2214_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2931_ (.I(_2228_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2932_ (.I(\mod.instr_2[14] ),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2933_ (.I(_2230_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2934_ (.I(_2197_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2935_ (.I(_2232_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2936_ (.A1(_2231_),
    .A2(_2227_),
    .A3(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2937_ (.I(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2938_ (.A1(\mod.registers.r4[15] ),
    .A2(_2229_),
    .B1(_2235_),
    .B2(\mod.registers.r1[15] ),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2939_ (.A1(_2217_),
    .A2(_2226_),
    .A3(_2236_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2940_ (.I(\mod.funct7[2] ),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2941_ (.I(\mod.instr_2[1] ),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2942_ (.I(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2943_ (.A1(_2238_),
    .A2(_2188_),
    .B(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2944_ (.A1(_2190_),
    .A2(_2237_),
    .B(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2945_ (.I(\mod.funct7[1] ),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2946_ (.I(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2947_ (.I(_2240_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2948_ (.I(_2245_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2949_ (.I(_2188_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2950_ (.A1(_2244_),
    .A2(_2246_),
    .A3(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2951_ (.A1(_2242_),
    .A2(_2248_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2952_ (.A1(_2186_),
    .A2(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2953_ (.I(\mod.funct3[2] ),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2954_ (.I(_2251_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2955_ (.I(_2252_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2956_ (.I(\mod.funct3[1] ),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2957_ (.A1(\mod.instr_2[2] ),
    .A2(_2127_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2958_ (.I(_2255_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2959_ (.A1(_2239_),
    .A2(_2188_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2960_ (.I(_2257_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2961_ (.I(_2258_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2962_ (.A1(_2256_),
    .A2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2963_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2964_ (.A1(_2253_),
    .A2(_2254_),
    .A3(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2965_ (.I(_2262_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2966_ (.I(_2263_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2967_ (.I(_2257_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2968_ (.I(_2265_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2969_ (.I(_2266_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2970_ (.I(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2971_ (.I(_2191_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2972_ (.I(_2269_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2973_ (.A1(_2124_),
    .A2(\mod.instr_2[0] ),
    .B(\mod.instr_2[1] ),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2974_ (.I(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2975_ (.A1(_2256_),
    .A2(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2976_ (.I(_2273_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2977_ (.I(_2274_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2978_ (.A1(_2238_),
    .A2(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2979_ (.I(_2276_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2980_ (.A1(_2270_),
    .A2(_2275_),
    .B(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2981_ (.A1(\mod.registers.r5[13] ),
    .A2(_2201_),
    .B1(_2210_),
    .B2(\mod.registers.r2[13] ),
    .C1(_2216_),
    .C2(\mod.registers.r6[13] ),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2982_ (.A1(\mod.registers.r7[13] ),
    .A2(_2220_),
    .B1(_2225_),
    .B2(\mod.registers.r3[13] ),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2983_ (.A1(\mod.registers.r4[13] ),
    .A2(_2229_),
    .B1(_2235_),
    .B2(\mod.registers.r1[13] ),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2984_ (.A1(_2279_),
    .A2(_2280_),
    .A3(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2985_ (.A1(_2189_),
    .A2(_2282_),
    .B(_2241_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2986_ (.A1(\mod.registers.r7[13] ),
    .A2(_2169_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2987_ (.A1(_2142_),
    .A2(_2163_),
    .A3(_2157_),
    .A4(\mod.registers.r1[13] ),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2988_ (.I(\mod.instr_2[11] ),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2989_ (.I(_2286_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2990_ (.I(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2991_ (.I(_2161_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2992_ (.I(_2289_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2993_ (.I(_2143_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2994_ (.I(_2291_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2995_ (.I(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2996_ (.A1(_2288_),
    .A2(_2290_),
    .A3(_2293_),
    .A4(\mod.registers.r5[13] ),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2997_ (.I(_2174_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2998_ (.I(_2295_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2999_ (.A1(_2288_),
    .A2(_2172_),
    .A3(_2296_),
    .A4(\mod.registers.r6[13] ),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3000_ (.A1(_2284_),
    .A2(_2285_),
    .A3(_2294_),
    .A4(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3001_ (.I(_2133_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3002_ (.I(_2299_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3003_ (.I(_2300_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3004_ (.A1(_2288_),
    .A2(_2163_),
    .A3(_2177_),
    .A4(\mod.registers.r4[13] ),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3005_ (.A1(_2142_),
    .A2(_2172_),
    .A3(_2177_),
    .A4(\mod.registers.r2[13] ),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3006_ (.A1(_2142_),
    .A2(\mod.registers.r3[13] ),
    .A3(_2146_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3007_ (.A1(_2301_),
    .A2(_2302_),
    .A3(_2303_),
    .A4(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3008_ (.A1(\mod.pc_2[13] ),
    .A2(_2136_),
    .B1(_2298_),
    .B2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3009_ (.I(_2306_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3010_ (.A1(_2268_),
    .A2(_2278_),
    .B(_2283_),
    .C(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3011_ (.I(_2259_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3012_ (.A1(_2309_),
    .A2(_2278_),
    .B(_2283_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3013_ (.A1(_2307_),
    .A2(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3014_ (.A1(_2307_),
    .A2(_2310_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3015_ (.A1(_2311_),
    .A2(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3016_ (.I(\mod.registers.r1[12] ),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3017_ (.I(_2160_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3018_ (.A1(_2140_),
    .A2(_2315_),
    .A3(_2155_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3019_ (.I(_2316_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3020_ (.I(_2166_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3021_ (.I(_2160_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3022_ (.A1(_2318_),
    .A2(_2319_),
    .A3(_2292_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3023_ (.I(\mod.registers.r5[12] ),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3024_ (.A1(_2314_),
    .A2(_2317_),
    .B1(_2320_),
    .B2(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3025_ (.I(\mod.registers.r6[12] ),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3026_ (.I(_2286_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3027_ (.I(_2151_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3028_ (.I(_2325_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3029_ (.A1(_2324_),
    .A2(_2326_),
    .A3(_2295_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3030_ (.A1(\mod.registers.r7[12] ),
    .A2(_2169_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3031_ (.A1(_2323_),
    .A2(_2327_),
    .B(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3032_ (.I(_2139_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3033_ (.I(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3034_ (.I(_2326_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3035_ (.A1(_2331_),
    .A2(_2332_),
    .A3(_2296_),
    .A4(\mod.registers.r2[12] ),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3036_ (.A1(_2331_),
    .A2(\mod.registers.r3[12] ),
    .A3(_2146_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3037_ (.A1(_2288_),
    .A2(_2290_),
    .A3(_2296_),
    .A4(\mod.registers.r4[12] ),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3038_ (.A1(_2135_),
    .A2(_2333_),
    .A3(_2334_),
    .A4(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3039_ (.A1(_2322_),
    .A2(_2329_),
    .A3(_2336_),
    .B1(_2301_),
    .B2(\mod.pc_2[12] ),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3040_ (.I(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3041_ (.I(_2132_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3042_ (.A1(\mod.funct7[2] ),
    .A2(_2239_),
    .A3(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3043_ (.A1(_2257_),
    .A2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3044_ (.I(_2341_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3045_ (.A1(\mod.registers.r4[12] ),
    .A2(_2229_),
    .B1(_2225_),
    .B2(\mod.registers.r3[12] ),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3046_ (.A1(\mod.registers.r5[12] ),
    .A2(_2201_),
    .B1(_2210_),
    .B2(\mod.registers.r2[12] ),
    .C1(_2216_),
    .C2(\mod.registers.r6[12] ),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3047_ (.A1(\mod.registers.r7[12] ),
    .A2(_2220_),
    .B1(_2235_),
    .B2(\mod.registers.r1[12] ),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3048_ (.A1(_2343_),
    .A2(_2344_),
    .A3(_2345_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3049_ (.A1(_2189_),
    .A2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3050_ (.I(_2205_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3051_ (.A1(_2348_),
    .A2(_2275_),
    .B(_2276_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3052_ (.A1(_2342_),
    .A2(_2347_),
    .B1(_2349_),
    .B2(_2309_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3053_ (.I(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3054_ (.A1(_2338_),
    .A2(_2351_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3055_ (.I(_2352_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3056_ (.A1(_2313_),
    .A2(_2353_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3057_ (.I(_2271_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3058_ (.I(_2355_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3059_ (.I(_2198_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3060_ (.A1(_2193_),
    .A2(_2196_),
    .A3(_2357_),
    .A4(\mod.registers.r2[0] ),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3061_ (.I(_2222_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3062_ (.A1(_2221_),
    .A2(\mod.registers.r3[0] ),
    .A3(_2359_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3063_ (.I(_2230_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3064_ (.I(_2212_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3065_ (.A1(_2361_),
    .A2(_2362_),
    .A3(_2199_),
    .A4(\mod.registers.r4[0] ),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3066_ (.A1(_2358_),
    .A2(_2360_),
    .A3(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3067_ (.I(_2218_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3068_ (.A1(\mod.registers.r7[0] ),
    .A2(_2365_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3069_ (.I(_2230_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3070_ (.A1(_2367_),
    .A2(_2213_),
    .A3(_2208_),
    .A4(\mod.registers.r5[0] ),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3071_ (.A1(_2367_),
    .A2(_2196_),
    .A3(_2357_),
    .A4(\mod.registers.r6[0] ),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3072_ (.A1(_2193_),
    .A2(_2362_),
    .A3(_2214_),
    .A4(\mod.registers.r1[0] ),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3073_ (.A1(_2366_),
    .A2(_2368_),
    .A3(_2369_),
    .A4(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3074_ (.I(\mod.instr_2[3] ),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3075_ (.A1(\mod.funct3[2] ),
    .A2(_2255_),
    .B(_2132_),
    .C(_2239_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3076_ (.I(_2373_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3077_ (.A1(_2124_),
    .A2(_2127_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3078_ (.A1(_2251_),
    .A2(_2375_),
    .B(_2272_),
    .C(_2208_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3079_ (.I(_2272_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3080_ (.A1(_2372_),
    .A2(_2374_),
    .B(_2376_),
    .C(_2377_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3081_ (.A1(_2356_),
    .A2(_2364_),
    .A3(_2371_),
    .B(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3082_ (.A1(_2266_),
    .A2(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3083_ (.I(\mod.registers.r3[0] ),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3084_ (.A1(_2140_),
    .A2(_2145_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3085_ (.I(_2166_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3086_ (.A1(_2383_),
    .A2(_2315_),
    .A3(_2175_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3087_ (.I(\mod.registers.r4[0] ),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3088_ (.A1(_2381_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3089_ (.I(\mod.registers.r1[0] ),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3090_ (.A1(\mod.registers.r7[0] ),
    .A2(_2168_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3091_ (.A1(_2387_),
    .A2(_2316_),
    .B(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3092_ (.I(_2299_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3093_ (.I(_2383_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3094_ (.I(_2291_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3095_ (.A1(_2391_),
    .A2(_2162_),
    .A3(_2392_),
    .A4(\mod.registers.r5[0] ),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3096_ (.I(_2325_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3097_ (.I(_2173_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3098_ (.I(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3099_ (.A1(_2391_),
    .A2(_2394_),
    .A3(_2396_),
    .A4(\mod.registers.r6[0] ),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3100_ (.A1(_2141_),
    .A2(_2171_),
    .A3(_2396_),
    .A4(\mod.registers.r2[0] ),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3101_ (.A1(_2390_),
    .A2(_2393_),
    .A3(_2397_),
    .A4(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3102_ (.I(\mod.pc_2[0] ),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3103_ (.A1(_2400_),
    .A2(_2265_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3104_ (.A1(_2386_),
    .A2(_2389_),
    .A3(_2399_),
    .B(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3105_ (.I(_2402_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3106_ (.I(_2355_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3107_ (.I(\mod.registers.r2[1] ),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3108_ (.A1(_2191_),
    .A2(_2195_),
    .A3(_2198_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3109_ (.I(_2406_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3110_ (.I(_2192_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3111_ (.A1(_2408_),
    .A2(\mod.registers.r3[1] ),
    .A3(_2223_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3112_ (.I(_2230_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3113_ (.A1(_2410_),
    .A2(_2362_),
    .A3(_2199_),
    .A4(\mod.registers.r4[1] ),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3114_ (.A1(_2405_),
    .A2(_2407_),
    .B(_2409_),
    .C(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3115_ (.I(_2218_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3116_ (.A1(\mod.registers.r7[1] ),
    .A2(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3117_ (.I(_2212_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3118_ (.A1(_2410_),
    .A2(_2415_),
    .A3(_2214_),
    .A4(\mod.registers.r5[1] ),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3119_ (.A1(_2410_),
    .A2(_2227_),
    .A3(_2233_),
    .A4(\mod.registers.r6[1] ),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3120_ (.I(_2207_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3121_ (.A1(_2408_),
    .A2(_2415_),
    .A3(_2418_),
    .A4(\mod.registers.r1[1] ),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3122_ (.A1(_2414_),
    .A2(_2416_),
    .A3(_2417_),
    .A4(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3123_ (.I(\mod.instr_2[4] ),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3124_ (.I(_2195_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3125_ (.A1(_2251_),
    .A2(_2375_),
    .B(_2272_),
    .C(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3126_ (.A1(_2421_),
    .A2(_2374_),
    .B(_2423_),
    .C(_2377_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3127_ (.A1(_2404_),
    .A2(_2412_),
    .A3(_2420_),
    .B(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3128_ (.I(_2174_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3129_ (.A1(_2324_),
    .A2(_2289_),
    .A3(_2426_),
    .A4(\mod.registers.r4[1] ),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3130_ (.I(_2139_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3131_ (.I(_2144_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3132_ (.A1(_2428_),
    .A2(\mod.registers.r3[1] ),
    .A3(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3133_ (.A1(_2427_),
    .A2(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3134_ (.I(_2133_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3135_ (.A1(_2330_),
    .A2(_2289_),
    .A3(_2292_),
    .A4(\mod.registers.r1[1] ),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3136_ (.A1(_2432_),
    .A2(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3137_ (.I(_2151_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3138_ (.A1(_2148_),
    .A2(_2435_),
    .A3(_2426_),
    .A4(\mod.registers.r2[1] ),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3139_ (.I(_2167_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3140_ (.A1(\mod.registers.r7[1] ),
    .A2(_2437_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3141_ (.I(_2174_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3142_ (.A1(_2318_),
    .A2(_2435_),
    .A3(_2439_),
    .A4(\mod.registers.r6[1] ),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3143_ (.I(_2291_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3144_ (.A1(_2318_),
    .A2(_2319_),
    .A3(_2441_),
    .A4(\mod.registers.r5[1] ),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3145_ (.A1(_2436_),
    .A2(_2438_),
    .A3(_2440_),
    .A4(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3146_ (.I(\mod.pc_2[1] ),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3147_ (.I(_2257_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3148_ (.A1(_2444_),
    .A2(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3149_ (.A1(_2431_),
    .A2(_2434_),
    .A3(_2443_),
    .B(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3150_ (.I(_2447_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3151_ (.A1(_2259_),
    .A2(_2425_),
    .B(_2448_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3152_ (.A1(\mod.registers.r4[1] ),
    .A2(_2228_),
    .B1(_2209_),
    .B2(\mod.registers.r2[1] ),
    .C1(_2224_),
    .C2(\mod.registers.r3[1] ),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3153_ (.A1(_2414_),
    .A2(_2416_),
    .A3(_2417_),
    .A4(_2419_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3154_ (.A1(_2450_),
    .A2(_2451_),
    .B(_2131_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3155_ (.A1(_2421_),
    .A2(_2374_),
    .B(_2423_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3156_ (.A1(_2356_),
    .A2(_2453_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3157_ (.I(_2445_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3158_ (.A1(_2427_),
    .A2(_2430_),
    .A3(_2438_),
    .A4(_2433_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3159_ (.A1(_2300_),
    .A2(_2436_),
    .A3(_2440_),
    .A4(_2442_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3160_ (.A1(_2444_),
    .A2(_2455_),
    .B1(_2456_),
    .B2(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3161_ (.A1(_2452_),
    .A2(_2454_),
    .B(_2458_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3162_ (.A1(_2380_),
    .A2(_2403_),
    .B1(_2449_),
    .B2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3163_ (.I(_2265_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3164_ (.A1(_2461_),
    .A2(_2425_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3165_ (.A1(_2462_),
    .A2(_2448_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3166_ (.I0(\mod.instr_2[5] ),
    .I1(_2361_),
    .S(_2373_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3167_ (.I(\mod.registers.r5[2] ),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3168_ (.A1(_2202_),
    .A2(_2204_),
    .A3(_2206_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3169_ (.I(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3170_ (.I(\mod.registers.r2[2] ),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3171_ (.I(_2202_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3172_ (.I(_2194_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3173_ (.A1(_2469_),
    .A2(_2470_),
    .A3(_2232_),
    .A4(\mod.registers.r6[2] ),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3174_ (.A1(_2465_),
    .A2(_2467_),
    .B1(_2406_),
    .B2(_2468_),
    .C(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3175_ (.I(_2191_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3176_ (.I(_2204_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3177_ (.I(_2207_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3178_ (.A1(_2473_),
    .A2(_2474_),
    .A3(_2475_),
    .A4(\mod.registers.r1[2] ),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3179_ (.A1(_2473_),
    .A2(\mod.registers.r3[2] ),
    .A3(_2222_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3180_ (.A1(_2469_),
    .A2(_2474_),
    .A3(_2232_),
    .A4(\mod.registers.r4[2] ),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3181_ (.A1(\mod.registers.r7[2] ),
    .A2(_2218_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3182_ (.A1(_2476_),
    .A2(_2477_),
    .A3(_2478_),
    .A4(_2479_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _3183_ (.A1(_2240_),
    .A2(_2339_),
    .A3(_2464_),
    .B1(_2472_),
    .B2(_2480_),
    .B3(_2355_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3184_ (.A1(_2258_),
    .A2(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3185_ (.I(_2432_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3186_ (.I(_2161_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3187_ (.A1(_2428_),
    .A2(_2484_),
    .A3(_2292_),
    .A4(\mod.registers.r1[2] ),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3188_ (.A1(_2428_),
    .A2(\mod.registers.r3[2] ),
    .A3(_2429_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3189_ (.A1(\mod.registers.r7[2] ),
    .A2(_2437_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3190_ (.I(_2286_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3191_ (.A1(_2488_),
    .A2(_2289_),
    .A3(_2295_),
    .A4(\mod.registers.r4[2] ),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3192_ (.A1(_2485_),
    .A2(_2486_),
    .A3(_2487_),
    .A4(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3193_ (.A1(_2488_),
    .A2(_2484_),
    .A3(_2392_),
    .A4(\mod.registers.r5[2] ),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3194_ (.A1(_2488_),
    .A2(_2326_),
    .A3(_2295_),
    .A4(\mod.registers.r6[2] ),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3195_ (.I(_2138_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3196_ (.I(_2493_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3197_ (.I(_2395_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3198_ (.A1(_2494_),
    .A2(_2326_),
    .A3(_2495_),
    .A4(\mod.registers.r2[2] ),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3199_ (.A1(_2134_),
    .A2(_2491_),
    .A3(_2492_),
    .A4(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3200_ (.A1(\mod.pc_2[2] ),
    .A2(_2483_),
    .B1(_2490_),
    .B2(_2497_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3201_ (.A1(_2482_),
    .A2(_2498_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3202_ (.A1(_2460_),
    .A2(_2463_),
    .B(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3203_ (.I(\mod.funct7[0] ),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3204_ (.A1(\mod.registers.r7[3] ),
    .A2(_2219_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3205_ (.A1(\mod.registers.r1[3] ),
    .A2(_2234_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3206_ (.A1(\mod.registers.r5[3] ),
    .A2(_2200_),
    .B1(_2209_),
    .B2(\mod.registers.r2[3] ),
    .C1(_2215_),
    .C2(\mod.registers.r6[3] ),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3207_ (.A1(\mod.registers.r4[3] ),
    .A2(_2228_),
    .B1(_2224_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3208_ (.A1(_2502_),
    .A2(_2503_),
    .A3(_2504_),
    .A4(_2505_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3209_ (.A1(_2501_),
    .A2(_2189_),
    .B1(_2506_),
    .B2(_2187_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3210_ (.I(\mod.registers.r3[3] ),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3211_ (.I(_2382_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3212_ (.I(_2384_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3213_ (.I(\mod.registers.r4[3] ),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3214_ (.A1(_2508_),
    .A2(_2509_),
    .B1(_2510_),
    .B2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3215_ (.I(\mod.registers.r1[3] ),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3216_ (.A1(_2513_),
    .A2(_2317_),
    .B(_2483_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3217_ (.I(_2167_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3218_ (.A1(\mod.registers.r7[3] ),
    .A2(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3219_ (.I(_2324_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3220_ (.A1(_2517_),
    .A2(_2290_),
    .A3(_2293_),
    .A4(\mod.registers.r5[3] ),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3221_ (.I(_2439_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3222_ (.A1(_2517_),
    .A2(_2153_),
    .A3(_2519_),
    .A4(\mod.registers.r6[3] ),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3223_ (.A1(_2331_),
    .A2(_2332_),
    .A3(_2519_),
    .A4(\mod.registers.r2[3] ),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3224_ (.A1(_2516_),
    .A2(_2518_),
    .A3(_2520_),
    .A4(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3225_ (.I(\mod.pc_2[3] ),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3226_ (.A1(_2523_),
    .A2(_2258_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3227_ (.A1(_2512_),
    .A2(_2514_),
    .A3(_2522_),
    .B(_2524_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3228_ (.A1(_2507_),
    .A2(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3229_ (.I(_2498_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3230_ (.A1(_2482_),
    .A2(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3231_ (.A1(_2526_),
    .A2(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3232_ (.I(\mod.registers.r5[7] ),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3233_ (.I(_2197_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3234_ (.A1(_2469_),
    .A2(_2470_),
    .A3(_2531_),
    .A4(\mod.registers.r6[7] ),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3235_ (.A1(_2203_),
    .A2(_2205_),
    .A3(_2531_),
    .A4(\mod.registers.r4[7] ),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3236_ (.A1(_2530_),
    .A2(_2467_),
    .B(_2532_),
    .C(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3237_ (.A1(\mod.registers.r7[7] ),
    .A2(_2365_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3238_ (.I(_2198_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3239_ (.A1(_2269_),
    .A2(_2422_),
    .A3(_2536_),
    .A4(\mod.registers.r2[7] ),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3240_ (.A1(_2211_),
    .A2(\mod.registers.r3[7] ),
    .A3(_2359_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3241_ (.A1(_2211_),
    .A2(_2205_),
    .A3(_2475_),
    .A4(\mod.registers.r1[7] ),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3242_ (.A1(_2535_),
    .A2(_2537_),
    .A3(_2538_),
    .A4(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3243_ (.A1(_2377_),
    .A2(_2534_),
    .A3(_2540_),
    .B(_2341_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3244_ (.I(_2273_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3245_ (.A1(_2251_),
    .A2(_2273_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3246_ (.A1(_2542_),
    .A2(_2464_),
    .B(_2543_),
    .C(_2445_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3247_ (.A1(\mod.registers.r7[7] ),
    .A2(_2437_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3248_ (.I(_2160_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3249_ (.A1(_2148_),
    .A2(_2546_),
    .A3(_2441_),
    .A4(\mod.registers.r1[7] ),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3250_ (.A1(_2179_),
    .A2(_2319_),
    .A3(_2441_),
    .A4(\mod.registers.r5[7] ),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3251_ (.A1(_2318_),
    .A2(_2435_),
    .A3(_2439_),
    .A4(\mod.registers.r6[7] ),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3252_ (.A1(_2545_),
    .A2(_2547_),
    .A3(_2548_),
    .A4(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3253_ (.A1(_2324_),
    .A2(_2319_),
    .A3(_2426_),
    .A4(\mod.registers.r4[7] ),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3254_ (.A1(_2330_),
    .A2(_2435_),
    .A3(_2426_),
    .A4(\mod.registers.r2[7] ),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3255_ (.A1(_2330_),
    .A2(\mod.registers.r3[7] ),
    .A3(_2145_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3256_ (.A1(_2432_),
    .A2(_0264_),
    .A3(_0265_),
    .A4(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3257_ (.A1(\mod.pc_2[7] ),
    .A2(_2390_),
    .B1(_2550_),
    .B2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3258_ (.A1(_2541_),
    .A2(_2544_),
    .B(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3259_ (.A1(_0268_),
    .A2(_2541_),
    .A3(_2544_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3260_ (.A1(_0269_),
    .A2(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3261_ (.I(\mod.registers.r4[6] ),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3262_ (.A1(_0272_),
    .A2(_2384_),
    .B(_2299_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3263_ (.A1(_2179_),
    .A2(_2546_),
    .A3(_2441_),
    .A4(\mod.registers.r5[6] ),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3264_ (.A1(_2179_),
    .A2(_2152_),
    .A3(_2439_),
    .A4(\mod.registers.r6[6] ),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3265_ (.A1(\mod.registers.r7[6] ),
    .A2(_2437_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3266_ (.A1(_2148_),
    .A2(_2546_),
    .A3(_2155_),
    .A4(\mod.registers.r1[6] ),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3267_ (.A1(_0274_),
    .A2(_0275_),
    .A3(_0276_),
    .A4(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3268_ (.I(\mod.registers.r3[6] ),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3269_ (.A1(_2493_),
    .A2(_2152_),
    .A3(_2175_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3270_ (.I(\mod.registers.r2[6] ),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3271_ (.A1(_0279_),
    .A2(_2382_),
    .B1(_0280_),
    .B2(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3272_ (.A1(_0273_),
    .A2(_0278_),
    .A3(_0282_),
    .B1(_2134_),
    .B2(\mod.pc_2[6] ),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3273_ (.I(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3274_ (.I(\mod.registers.r5[6] ),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3275_ (.A1(_2269_),
    .A2(_2474_),
    .A3(_2475_),
    .A4(\mod.registers.r1[6] ),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3276_ (.A1(\mod.registers.r7[6] ),
    .A2(_2365_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3277_ (.A1(_0285_),
    .A2(_2467_),
    .B(_0286_),
    .C(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3278_ (.A1(_2367_),
    .A2(_2213_),
    .A3(_2536_),
    .A4(\mod.registers.r4[6] ),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3279_ (.A1(_2211_),
    .A2(\mod.registers.r3[6] ),
    .A3(_2359_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3280_ (.A1(_2269_),
    .A2(_2422_),
    .A3(_2536_),
    .A4(\mod.registers.r2[6] ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3281_ (.A1(_2367_),
    .A2(_2196_),
    .A3(_2357_),
    .A4(\mod.registers.r6[6] ),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3282_ (.A1(_0289_),
    .A2(_0290_),
    .A3(_0291_),
    .A4(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3283_ (.A1(_2377_),
    .A2(_0288_),
    .A3(_0293_),
    .B(_2341_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3284_ (.A1(_2256_),
    .A2(_2271_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3285_ (.A1(\mod.funct3[1] ),
    .A2(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3286_ (.A1(_2542_),
    .A2(_2453_),
    .B(_0296_),
    .C(_2445_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3287_ (.A1(_0294_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3288_ (.A1(_0284_),
    .A2(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3289_ (.I(\mod.registers.r5[5] ),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3290_ (.I(_2466_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3291_ (.I(\mod.registers.r2[5] ),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3292_ (.A1(_2361_),
    .A2(_2227_),
    .A3(_2199_),
    .A4(\mod.registers.r6[5] ),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3293_ (.A1(_0300_),
    .A2(_0301_),
    .B1(_2407_),
    .B2(_0302_),
    .C(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3294_ (.A1(\mod.registers.r7[5] ),
    .A2(_2413_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3295_ (.A1(_2408_),
    .A2(\mod.registers.r3[5] ),
    .A3(_2223_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3296_ (.A1(_2408_),
    .A2(_2415_),
    .A3(_2418_),
    .A4(\mod.registers.r1[5] ),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3297_ (.A1(_2410_),
    .A2(_2415_),
    .A3(_2233_),
    .A4(\mod.registers.r4[5] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3298_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0307_),
    .A4(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3299_ (.A1(_2404_),
    .A2(_0304_),
    .A3(_0309_),
    .B(_2341_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3300_ (.A1(_2372_),
    .A2(_2374_),
    .B(_2376_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3301_ (.I(\mod.funct3[0] ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3302_ (.A1(_0312_),
    .A2(_2542_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3303_ (.A1(_2542_),
    .A2(_0311_),
    .B(_0313_),
    .C(_2265_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3304_ (.A1(_2286_),
    .A2(_2161_),
    .A3(_2395_),
    .A4(\mod.registers.r4[5] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3305_ (.A1(\mod.registers.r7[5] ),
    .A2(_2167_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3306_ (.A1(_2493_),
    .A2(_2325_),
    .A3(_2395_),
    .A4(\mod.registers.r2[5] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3307_ (.A1(_2493_),
    .A2(\mod.registers.r3[5] ),
    .A3(_2145_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3308_ (.A1(_0315_),
    .A2(_0316_),
    .A3(_0317_),
    .A4(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3309_ (.A1(_2383_),
    .A2(_2325_),
    .A3(_2175_),
    .A4(\mod.registers.r6[5] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3310_ (.A1(_2383_),
    .A2(_2315_),
    .A3(_2291_),
    .A4(\mod.registers.r5[5] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3311_ (.A1(_2140_),
    .A2(_2315_),
    .A3(_2155_),
    .A4(\mod.registers.r1[5] ),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3312_ (.A1(_2299_),
    .A2(_0320_),
    .A3(_0321_),
    .A4(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3313_ (.A1(\mod.pc_2[5] ),
    .A2(_2432_),
    .B1(_0319_),
    .B2(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3314_ (.I(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3315_ (.A1(_0310_),
    .A2(_0314_),
    .B(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3316_ (.A1(_0324_),
    .A2(_0310_),
    .A3(_0314_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3317_ (.A1(_0326_),
    .A2(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3318_ (.A1(_2494_),
    .A2(_2394_),
    .A3(_2495_),
    .A4(\mod.registers.r2[4] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3319_ (.A1(_2428_),
    .A2(_2484_),
    .A3(_2392_),
    .A4(\mod.registers.r1[4] ),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3320_ (.A1(\mod.registers.r7[4] ),
    .A2(_2168_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3321_ (.A1(_2287_),
    .A2(_2162_),
    .A3(_2495_),
    .A4(\mod.registers.r4[4] ),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3322_ (.A1(_0329_),
    .A2(_0330_),
    .A3(_0331_),
    .A4(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3323_ (.A1(_2287_),
    .A2(_2394_),
    .A3(_2396_),
    .A4(\mod.registers.r6[4] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3324_ (.A1(_2141_),
    .A2(\mod.registers.r3[4] ),
    .A3(_2429_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3325_ (.A1(_2287_),
    .A2(_2162_),
    .A3(_2392_),
    .A4(\mod.registers.r5[4] ),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3326_ (.A1(_2390_),
    .A2(_0334_),
    .A3(_0335_),
    .A4(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3327_ (.A1(\mod.pc_2[4] ),
    .A2(_2135_),
    .B1(_0333_),
    .B2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3328_ (.I(\mod.registers.r5[4] ),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3329_ (.I(\mod.registers.r2[4] ),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3330_ (.A1(_2203_),
    .A2(_2422_),
    .A3(_2536_),
    .A4(\mod.registers.r6[4] ),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3331_ (.A1(_0339_),
    .A2(_2467_),
    .B1(_2406_),
    .B2(_0340_),
    .C(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3332_ (.A1(_2221_),
    .A2(\mod.registers.r3[4] ),
    .A3(_2359_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3333_ (.A1(_2193_),
    .A2(_2213_),
    .A3(_2208_),
    .A4(\mod.registers.r1[4] ),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3334_ (.A1(_2361_),
    .A2(_2362_),
    .A3(_2357_),
    .A4(\mod.registers.r4[4] ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3335_ (.A1(\mod.registers.r7[4] ),
    .A2(_2365_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3336_ (.A1(_0343_),
    .A2(_0344_),
    .A3(_0345_),
    .A4(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _3337_ (.A1(\mod.funct7[1] ),
    .A2(_2240_),
    .A3(_2339_),
    .B1(_2404_),
    .B2(_0342_),
    .B3(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3338_ (.A1(_2461_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3339_ (.A1(_0333_),
    .A2(_0337_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3340_ (.A1(_2266_),
    .A2(_0350_),
    .A3(_0348_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3341_ (.A1(_0338_),
    .A2(_0349_),
    .B(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3342_ (.A1(_0271_),
    .A2(_0299_),
    .A3(_0328_),
    .A4(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3343_ (.I(_2525_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3344_ (.A1(_2507_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3345_ (.A1(_2500_),
    .A2(_2529_),
    .B(_0353_),
    .C(_0355_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3346_ (.I(_0271_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3347_ (.A1(_0284_),
    .A2(_0294_),
    .A3(_0297_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3348_ (.A1(_2550_),
    .A2(_0267_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3349_ (.A1(\mod.pc_2[7] ),
    .A2(_2301_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3350_ (.A1(_0359_),
    .A2(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3351_ (.A1(_0361_),
    .A2(_2541_),
    .A3(_2544_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3352_ (.A1(_0357_),
    .A2(_0358_),
    .B(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3353_ (.A1(_0319_),
    .A2(_0323_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3354_ (.A1(\mod.pc_2[5] ),
    .A2(_2301_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3355_ (.A1(_0364_),
    .A2(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3356_ (.A1(_0366_),
    .A2(_0310_),
    .A3(_0314_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3357_ (.I(_2355_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3358_ (.A1(_0342_),
    .A2(_0347_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3359_ (.A1(_2243_),
    .A2(_0368_),
    .B1(_0369_),
    .B2(_2246_),
    .C(_0338_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3360_ (.A1(_0326_),
    .A2(_0327_),
    .B(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3361_ (.A1(_0367_),
    .A2(_0371_),
    .B(_0357_),
    .C(_0299_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3362_ (.A1(_0363_),
    .A2(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3363_ (.A1(\mod.registers.r7[9] ),
    .A2(_2515_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3364_ (.I(_2546_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3365_ (.A1(_2149_),
    .A2(_0375_),
    .A3(_2156_),
    .A4(\mod.registers.r1[9] ),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3366_ (.A1(_2391_),
    .A2(_2171_),
    .A3(_2176_),
    .A4(\mod.registers.r6[9] ),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3367_ (.A1(_2180_),
    .A2(_0375_),
    .A3(_2156_),
    .A4(\mod.registers.r5[9] ),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3368_ (.A1(_0374_),
    .A2(_0376_),
    .A3(_0377_),
    .A4(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3369_ (.A1(_2149_),
    .A2(_2153_),
    .A3(_2176_),
    .A4(\mod.registers.r2[9] ),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3370_ (.A1(_2149_),
    .A2(\mod.registers.r3[9] ),
    .A3(_2146_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3371_ (.A1(_2180_),
    .A2(_0375_),
    .A3(_2519_),
    .A4(\mod.registers.r4[9] ),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3372_ (.A1(_2300_),
    .A2(_0380_),
    .A3(_0381_),
    .A4(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3373_ (.A1(_0379_),
    .A2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3374_ (.A1(\mod.pc_2[9] ),
    .A2(_2135_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3375_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3376_ (.I(\mod.registers.r5[9] ),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3377_ (.I(\mod.registers.r2[9] ),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3378_ (.I(_2470_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3379_ (.I(_2232_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3380_ (.A1(_2231_),
    .A2(_0389_),
    .A3(_0390_),
    .A4(\mod.registers.r6[9] ),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3381_ (.A1(_0387_),
    .A2(_0301_),
    .B1(_2407_),
    .B2(_0388_),
    .C(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3382_ (.I(_2473_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3383_ (.I(_2222_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3384_ (.A1(_0393_),
    .A2(\mod.registers.r3[9] ),
    .A3(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3385_ (.A1(\mod.registers.r7[9] ),
    .A2(_2219_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3386_ (.I(_2469_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3387_ (.I(_2212_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3388_ (.A1(_0397_),
    .A2(_0398_),
    .A3(_0390_),
    .A4(\mod.registers.r4[9] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3389_ (.I(_2474_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3390_ (.I(_2475_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3391_ (.A1(_0393_),
    .A2(_0400_),
    .A3(_0401_),
    .A4(\mod.registers.r1[9] ),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3392_ (.A1(_0395_),
    .A2(_0396_),
    .A3(_0399_),
    .A4(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3393_ (.A1(_2356_),
    .A2(_0392_),
    .A3(_0403_),
    .B(_2342_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3394_ (.I0(\mod.funct7[1] ),
    .I1(_2332_),
    .S(_2274_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3395_ (.A1(_2266_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3396_ (.A1(_0404_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3397_ (.A1(_0386_),
    .A2(_0407_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3398_ (.I(\mod.pc_2[11] ),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3399_ (.A1(\mod.registers.r7[11] ),
    .A2(_2515_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3400_ (.A1(_2180_),
    .A2(_2153_),
    .A3(_2519_),
    .A4(\mod.registers.r6[11] ),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3401_ (.A1(_2517_),
    .A2(_2290_),
    .A3(_2293_),
    .A4(\mod.registers.r5[11] ),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3402_ (.A1(_2331_),
    .A2(_2332_),
    .A3(_2296_),
    .A4(\mod.registers.r2[11] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3403_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0412_),
    .A4(_0413_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3404_ (.I(\mod.registers.r4[11] ),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3405_ (.A1(_0415_),
    .A2(_2510_),
    .B(_2483_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3406_ (.I(\mod.registers.r3[11] ),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3407_ (.I(\mod.registers.r1[11] ),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3408_ (.A1(_0417_),
    .A2(_2509_),
    .B1(_2317_),
    .B2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3409_ (.A1(_0416_),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3410_ (.A1(_0409_),
    .A2(_2461_),
    .B1(_0414_),
    .B2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3411_ (.I(_2531_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3412_ (.I(_2203_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3413_ (.A1(_0423_),
    .A2(_2348_),
    .A3(_0422_),
    .A4(\mod.registers.r4[11] ),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3414_ (.A1(_2270_),
    .A2(\mod.registers.r3[11] ),
    .A3(_0394_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(\mod.registers.r7[11] ),
    .A2(_2219_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3416_ (.A1(_0424_),
    .A2(_0425_),
    .A3(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3417_ (.I(_2470_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3418_ (.I(_2531_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3419_ (.A1(_2270_),
    .A2(_0428_),
    .A3(_0429_),
    .A4(\mod.registers.r2[11] ),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3420_ (.A1(_0397_),
    .A2(_0428_),
    .A3(_0429_),
    .A4(\mod.registers.r6[11] ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3421_ (.A1(_0423_),
    .A2(_0400_),
    .A3(_0401_),
    .A4(\mod.registers.r5[11] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3422_ (.A1(_0393_),
    .A2(_0400_),
    .A3(_0401_),
    .A4(\mod.registers.r1[11] ),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3423_ (.A1(_0430_),
    .A2(_0431_),
    .A3(_0432_),
    .A4(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3424_ (.A1(_0368_),
    .A2(_0427_),
    .A3(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3425_ (.A1(_0422_),
    .A2(_2245_),
    .A3(_2247_),
    .B1(_2241_),
    .B2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3426_ (.A1(_0421_),
    .A2(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3427_ (.I(\mod.registers.r5[10] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3428_ (.A1(\mod.registers.r7[10] ),
    .A2(_2413_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3429_ (.I(_2473_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3430_ (.A1(_0440_),
    .A2(_0398_),
    .A3(_2418_),
    .A4(\mod.registers.r1[10] ),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3431_ (.A1(_0438_),
    .A2(_0301_),
    .B(_0439_),
    .C(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3432_ (.A1(_0397_),
    .A2(_0400_),
    .A3(_0429_),
    .A4(\mod.registers.r4[10] ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3433_ (.A1(_0393_),
    .A2(\mod.registers.r3[10] ),
    .A3(_0394_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3434_ (.A1(_0440_),
    .A2(_0389_),
    .A3(_0390_),
    .A4(\mod.registers.r2[10] ),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3435_ (.A1(_0397_),
    .A2(_0389_),
    .A3(_0429_),
    .A4(\mod.registers.r6[10] ),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3436_ (.A1(_0443_),
    .A2(_0444_),
    .A3(_0445_),
    .A4(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3437_ (.A1(_0368_),
    .A2(_0442_),
    .A3(_0447_),
    .B(_2342_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3438_ (.I0(\mod.funct7[2] ),
    .I1(_2517_),
    .S(_2274_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3439_ (.A1(_2455_),
    .A2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3440_ (.I(\mod.registers.r3[10] ),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3441_ (.A1(_0451_),
    .A2(_2509_),
    .B1(_2320_),
    .B2(_0438_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3442_ (.I(\mod.registers.r4[10] ),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3443_ (.I(\mod.registers.r2[10] ),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3444_ (.A1(_0453_),
    .A2(_2510_),
    .B1(_0280_),
    .B2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3445_ (.A1(_2391_),
    .A2(_2171_),
    .A3(_2176_),
    .A4(\mod.registers.r6[10] ),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3446_ (.A1(\mod.registers.r7[10] ),
    .A2(_2515_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3447_ (.A1(_2141_),
    .A2(_0375_),
    .A3(_2156_),
    .A4(\mod.registers.r1[10] ),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3448_ (.A1(_2300_),
    .A2(_0456_),
    .A3(_0457_),
    .A4(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3449_ (.A1(\mod.pc_2[10] ),
    .A2(_2390_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3450_ (.A1(_0452_),
    .A2(_0455_),
    .A3(_0459_),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3451_ (.A1(_0448_),
    .A2(_0450_),
    .B(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3452_ (.A1(_0461_),
    .A2(_0448_),
    .A3(_0450_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3453_ (.A1(_0462_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3454_ (.I(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3455_ (.I(\mod.registers.r1[8] ),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3456_ (.I(\mod.registers.r5[8] ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3457_ (.A1(_0466_),
    .A2(_2316_),
    .B1(_2320_),
    .B2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3458_ (.I(\mod.registers.r6[8] ),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3459_ (.A1(\mod.registers.r7[8] ),
    .A2(_2168_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3460_ (.A1(_0469_),
    .A2(_2327_),
    .B(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3461_ (.A1(_2494_),
    .A2(_2394_),
    .A3(_2396_),
    .A4(\mod.registers.r2[8] ),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3462_ (.A1(_2494_),
    .A2(\mod.registers.r3[8] ),
    .A3(_2429_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3463_ (.A1(_2488_),
    .A2(_2484_),
    .A3(_2495_),
    .A4(\mod.registers.r4[8] ),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3464_ (.A1(_2134_),
    .A2(_0472_),
    .A3(_0473_),
    .A4(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3465_ (.A1(_0468_),
    .A2(_0471_),
    .A3(_0475_),
    .B1(_2483_),
    .B2(\mod.pc_2[8] ),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3466_ (.I(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3467_ (.I(\mod.registers.r2[8] ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3468_ (.A1(\mod.registers.r7[8] ),
    .A2(_2413_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3469_ (.A1(_0467_),
    .A2(_0301_),
    .B1(_2407_),
    .B2(_0478_),
    .C(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3470_ (.A1(_2231_),
    .A2(_0389_),
    .A3(_0390_),
    .A4(\mod.registers.r6[8] ),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3471_ (.A1(_2231_),
    .A2(_0398_),
    .A3(_2233_),
    .A4(\mod.registers.r4[8] ),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3472_ (.A1(_0440_),
    .A2(\mod.registers.r3[8] ),
    .A3(_2223_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3473_ (.A1(_0440_),
    .A2(_0398_),
    .A3(_2418_),
    .A4(\mod.registers.r1[8] ),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3474_ (.A1(_0481_),
    .A2(_0482_),
    .A3(_0483_),
    .A4(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3475_ (.A1(_2356_),
    .A2(_0480_),
    .A3(_0485_),
    .B(_2342_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3476_ (.I0(\mod.funct7[0] ),
    .I1(_2293_),
    .S(_2274_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3477_ (.A1(_2455_),
    .A2(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3478_ (.A1(_0486_),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3479_ (.A1(_0477_),
    .A2(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3480_ (.A1(_0408_),
    .A2(_0437_),
    .A3(_0465_),
    .A4(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3481_ (.A1(_0356_),
    .A2(_0373_),
    .B(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3482_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0412_),
    .A4(_0413_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3483_ (.A1(_0409_),
    .A2(_2461_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3484_ (.A1(_0493_),
    .A2(_0416_),
    .A3(_0419_),
    .B(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3485_ (.A1(_0495_),
    .A2(_0436_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3486_ (.I(_0461_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3487_ (.A1(_0497_),
    .A2(_0448_),
    .A3(_0450_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3488_ (.I(_0436_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3489_ (.A1(_0495_),
    .A2(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3490_ (.A1(_0496_),
    .A2(_0498_),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3491_ (.A1(_0437_),
    .A2(_0464_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3492_ (.I(_0477_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3493_ (.A1(_0503_),
    .A2(_0486_),
    .A3(_0488_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3494_ (.A1(_0386_),
    .A2(_0404_),
    .A3(_0406_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3495_ (.A1(_0408_),
    .A2(_0504_),
    .B(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3496_ (.A1(_0502_),
    .A2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3497_ (.A1(_0501_),
    .A2(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3498_ (.A1(_2338_),
    .A2(_2350_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3499_ (.A1(_2338_),
    .A2(_2350_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3500_ (.A1(_0509_),
    .A2(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3501_ (.A1(_0492_),
    .A2(_0508_),
    .B(_0511_),
    .C(_2313_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3502_ (.A1(\mod.registers.r5[14] ),
    .A2(_2201_),
    .B1(_2210_),
    .B2(\mod.registers.r2[14] ),
    .C1(_2216_),
    .C2(\mod.registers.r6[14] ),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3503_ (.A1(\mod.registers.r4[14] ),
    .A2(_2229_),
    .B1(_2225_),
    .B2(\mod.registers.r3[14] ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3504_ (.A1(\mod.registers.r7[14] ),
    .A2(_2220_),
    .B1(_2235_),
    .B2(\mod.registers.r1[14] ),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3505_ (.A1(_0513_),
    .A2(_0514_),
    .A3(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3506_ (.A1(_2190_),
    .A2(_0516_),
    .B(_2340_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3507_ (.A1(_2137_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3508_ (.I(\mod.registers.r3[14] ),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3509_ (.I(\mod.registers.r6[14] ),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3510_ (.A1(_0519_),
    .A2(_2509_),
    .B1(_2327_),
    .B2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3511_ (.I(\mod.registers.r1[14] ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3512_ (.A1(\mod.registers.r7[14] ),
    .A2(_2169_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3513_ (.A1(_0522_),
    .A2(_2317_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3514_ (.I(\mod.registers.r4[14] ),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3515_ (.I(\mod.registers.r2[14] ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3516_ (.I(\mod.registers.r5[14] ),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _3517_ (.A1(_0525_),
    .A2(_2510_),
    .B1(_0280_),
    .B2(_0526_),
    .C1(_2320_),
    .C2(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3518_ (.A1(_0521_),
    .A2(_0524_),
    .A3(_0528_),
    .B(_2136_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3519_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3520_ (.I(_2275_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3521_ (.A1(_2501_),
    .A2(_0531_),
    .B(_2277_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3522_ (.A1(_2268_),
    .A2(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3523_ (.A1(_0518_),
    .A2(_0530_),
    .A3(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3524_ (.A1(_2190_),
    .A2(_0516_),
    .B(_0530_),
    .C(_2340_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3525_ (.I(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3526_ (.A1(_0534_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3527_ (.A1(_2308_),
    .A2(_2354_),
    .A3(_0512_),
    .B(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3528_ (.A1(_0517_),
    .A2(_0530_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3529_ (.I(_2185_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3530_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3531_ (.A1(_2137_),
    .A2(_0540_),
    .B(_2249_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3532_ (.A1(_0541_),
    .A2(_2242_),
    .B(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3533_ (.I(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3534_ (.A1(_0538_),
    .A2(_0539_),
    .B(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3535_ (.A1(_0544_),
    .A2(_0538_),
    .A3(_0539_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3536_ (.A1(_2264_),
    .A2(_0545_),
    .A3(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3537_ (.I(_2482_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3538_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3539_ (.I(_0549_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3540_ (.A1(_2452_),
    .A2(_2454_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3541_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3542_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3543_ (.I(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3544_ (.I(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3545_ (.A1(\mod.pc_2[9] ),
    .A2(_2136_),
    .B1(_0379_),
    .B2(_0383_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3546_ (.A1(_2358_),
    .A2(_2360_),
    .A3(_2363_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3547_ (.A1(_2366_),
    .A2(_2368_),
    .A3(_2369_),
    .A4(_2370_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3548_ (.A1(_0557_),
    .A2(_0558_),
    .B(_2131_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3549_ (.A1(_2404_),
    .A2(_0311_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3550_ (.A1(_0559_),
    .A2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3551_ (.I(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3552_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3553_ (.I(_0561_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3554_ (.I(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3555_ (.A1(_0565_),
    .A2(_0503_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3556_ (.A1(_0556_),
    .A2(_0563_),
    .B(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3557_ (.I(_2380_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3558_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3559_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3560_ (.A1(_0495_),
    .A2(_0569_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3561_ (.A1(_0497_),
    .A2(_0570_),
    .B(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3562_ (.A1(_0555_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3563_ (.A1(_0555_),
    .A2(_0567_),
    .B(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3564_ (.I(_0563_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(_0551_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3566_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3567_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3568_ (.I(_2379_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3569_ (.A1(_2137_),
    .A2(_2185_),
    .A3(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3570_ (.A1(_0530_),
    .A2(_0575_),
    .B(_0578_),
    .C(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3571_ (.I(_2462_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3572_ (.I(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3573_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3574_ (.I(_2337_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3575_ (.A1(_2307_),
    .A2(_0570_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_0585_),
    .A2(_0570_),
    .B(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3577_ (.A1(_0584_),
    .A2(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3578_ (.A1(_0581_),
    .A2(_0588_),
    .B(_0550_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3579_ (.A1(_2502_),
    .A2(_2503_),
    .A3(_2504_),
    .A4(_2505_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3580_ (.A1(\mod.funct7[0] ),
    .A2(_0368_),
    .B1(_0590_),
    .B2(_2245_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3581_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3583_ (.I(\mod.funct3[2] ),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3584_ (.I(\mod.funct3[1] ),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3585_ (.A1(\mod.funct3[0] ),
    .A2(_2260_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3586_ (.A1(_0594_),
    .A2(_0595_),
    .A3(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3587_ (.I(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3588_ (.A1(_0593_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3589_ (.A1(_0550_),
    .A2(_0574_),
    .B(_0589_),
    .C(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3590_ (.I(_2462_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3591_ (.I(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3592_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3593_ (.I(_0283_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3594_ (.A1(_0361_),
    .A2(_0565_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3595_ (.A1(_0604_),
    .A2(_0563_),
    .B(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3596_ (.I(\mod.pc_2[4] ),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3597_ (.I(_2455_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3598_ (.A1(_0607_),
    .A2(_0608_),
    .B(_0350_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3599_ (.A1(_0325_),
    .A2(_0562_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3600_ (.A1(_0563_),
    .A2(_0609_),
    .B(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_0603_),
    .A2(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3602_ (.A1(_0603_),
    .A2(_0606_),
    .B(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3603_ (.I(_0559_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3604_ (.I(_0560_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3605_ (.A1(_0614_),
    .A2(_0615_),
    .B(_2402_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3606_ (.A1(_2268_),
    .A2(_0579_),
    .B(_2448_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3607_ (.A1(_0616_),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(_2527_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3609_ (.A1(_0619_),
    .A2(_0568_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3610_ (.I(_2267_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3611_ (.I(_2525_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3612_ (.A1(_0621_),
    .A2(_0579_),
    .B(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3613_ (.A1(_0620_),
    .A2(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3614_ (.I0(_0618_),
    .I1(_0624_),
    .S(_0577_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3615_ (.I(_2482_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3616_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3617_ (.I0(_0613_),
    .I1(_0625_),
    .S(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_2507_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3619_ (.I(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3620_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3621_ (.I(_0598_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3622_ (.A1(_0631_),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3623_ (.I(_2507_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3624_ (.A1(_0634_),
    .A2(_0548_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3625_ (.I(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3626_ (.I(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3627_ (.A1(_0584_),
    .A2(_0580_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3628_ (.A1(\mod.funct3[2] ),
    .A2(_2245_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3629_ (.A1(_2243_),
    .A2(_2128_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3630_ (.A1(_2125_),
    .A2(_0639_),
    .A3(_0640_),
    .B1(_2187_),
    .B2(_2375_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3631_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3632_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3633_ (.A1(_0637_),
    .A2(_0638_),
    .B(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3634_ (.I(_2254_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3635_ (.A1(_2253_),
    .A2(_0645_),
    .A3(_0596_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3636_ (.A1(_0541_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3637_ (.I(_0594_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3638_ (.A1(_0595_),
    .A2(\mod.funct3[0] ),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3639_ (.A1(_0648_),
    .A2(_2261_),
    .A3(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3640_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3641_ (.I(_0312_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3642_ (.A1(_0595_),
    .A2(_2260_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3643_ (.A1(_2252_),
    .A2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3644_ (.A1(_0652_),
    .A2(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3645_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3646_ (.I(\mod.funct3[0] ),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3647_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3648_ (.A1(_0658_),
    .A2(_0654_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3649_ (.A1(_0541_),
    .A2(_2242_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3650_ (.I(_2256_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3651_ (.A1(_2252_),
    .A2(_0649_),
    .B(_2268_),
    .C(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3652_ (.I(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3653_ (.A1(_0542_),
    .A2(_0656_),
    .B1(_0659_),
    .B2(_0660_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3654_ (.A1(_0543_),
    .A2(_0651_),
    .B(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3655_ (.A1(_0628_),
    .A2(_0633_),
    .B1(_0644_),
    .B2(_0647_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3656_ (.A1(_0600_),
    .A2(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3657_ (.A1(_2125_),
    .A2(_0639_),
    .A3(_0640_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3658_ (.A1(_2246_),
    .A2(_0661_),
    .B(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3659_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3660_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3661_ (.A1(_0545_),
    .A2(_0546_),
    .A3(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(_0591_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3663_ (.A1(_0673_),
    .A2(_0354_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3664_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3665_ (.A1(_2259_),
    .A2(_2425_),
    .A3(_2447_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3666_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3667_ (.I(_2379_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3668_ (.A1(_2267_),
    .A2(_0678_),
    .A3(_2403_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3669_ (.A1(_0677_),
    .A2(_0679_),
    .B(_2449_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3670_ (.A1(_0673_),
    .A2(_0354_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3671_ (.A1(_2258_),
    .A2(_2481_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3672_ (.I(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3673_ (.A1(_0683_),
    .A2(_2527_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3674_ (.A1(_2499_),
    .A2(_0680_),
    .B(_0681_),
    .C(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3675_ (.I(_0299_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3676_ (.I(_0352_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3677_ (.A1(_0357_),
    .A2(_0686_),
    .A3(_0328_),
    .A4(_0687_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3678_ (.A1(_0675_),
    .A2(_0685_),
    .A3(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3679_ (.I(_0269_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3680_ (.I(_0284_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3681_ (.I(_0298_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3682_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3683_ (.A1(_0325_),
    .A2(_0310_),
    .A3(_0314_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3684_ (.A1(_0691_),
    .A2(_0298_),
    .B1(_0326_),
    .B2(_0351_),
    .C(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3685_ (.A1(_0693_),
    .A2(_0695_),
    .B(_0270_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3686_ (.A1(_0690_),
    .A2(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3687_ (.I(_0437_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3688_ (.A1(_0698_),
    .A2(_0465_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3689_ (.I(_0490_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3690_ (.A1(_0408_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3691_ (.A1(_0699_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3692_ (.A1(_0689_),
    .A2(_0697_),
    .B(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3693_ (.I(_0421_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3694_ (.A1(_0704_),
    .A2(_0499_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3695_ (.I(_0462_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3696_ (.A1(_0404_),
    .A2(_0406_),
    .B(_0556_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3697_ (.A1(_0486_),
    .A2(_0488_),
    .B(_0476_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3698_ (.A1(_0556_),
    .A2(_0404_),
    .A3(_0406_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3699_ (.A1(_0707_),
    .A2(_0708_),
    .B(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3700_ (.A1(_0463_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3701_ (.A1(_0704_),
    .A2(_0499_),
    .B(_0706_),
    .C(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3702_ (.A1(_0705_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_0511_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3704_ (.A1(_2313_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3705_ (.A1(_0703_),
    .A2(_0713_),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3706_ (.A1(_2312_),
    .A2(_0585_),
    .A3(_2351_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3707_ (.A1(_2311_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3708_ (.I(_0537_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3709_ (.A1(_0716_),
    .A2(_0718_),
    .B(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3710_ (.I(_0544_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3711_ (.A1(_0536_),
    .A2(_0720_),
    .B(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3712_ (.A1(_0675_),
    .A2(_0685_),
    .A3(_0688_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3713_ (.A1(_0690_),
    .A2(_0696_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3714_ (.A1(_0723_),
    .A2(_0724_),
    .B(_0701_),
    .C(_0699_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3715_ (.A1(_0705_),
    .A2(_0712_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3716_ (.I(_2313_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3717_ (.A1(_0725_),
    .A2(_0726_),
    .B(_0727_),
    .C(_0714_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3718_ (.A1(_2311_),
    .A2(_0717_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3719_ (.A1(_0728_),
    .A2(_0729_),
    .B(_0537_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3720_ (.A1(_0544_),
    .A2(_0535_),
    .A3(_0730_),
    .B(_0671_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3721_ (.A1(_0648_),
    .A2(_2254_),
    .A3(_0657_),
    .B(_2261_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3722_ (.I(_0732_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3723_ (.I(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3724_ (.A1(_0722_),
    .A2(_0731_),
    .B(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3725_ (.A1(_0547_),
    .A2(_0667_),
    .B1(_0672_),
    .B2(_0735_),
    .C(_0721_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3726_ (.I(_0658_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3727_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3728_ (.A1(_2250_),
    .A2(_0736_),
    .B(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3729_ (.A1(_0737_),
    .A2(_2250_),
    .A3(_0736_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3730_ (.A1(_0739_),
    .A2(_0740_),
    .B(_0645_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3731_ (.A1(_0547_),
    .A2(_0667_),
    .B1(_0672_),
    .B2(_0735_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3732_ (.I(_0643_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3733_ (.A1(_2452_),
    .A2(_2454_),
    .A3(_2458_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3734_ (.A1(_0744_),
    .A2(_0676_),
    .B(_0616_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3735_ (.A1(_0552_),
    .A2(_2458_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3736_ (.A1(_0682_),
    .A2(_2498_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3737_ (.A1(_0745_),
    .A2(_0746_),
    .B(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3738_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3739_ (.A1(_2526_),
    .A2(_2528_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3740_ (.I(_0357_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3741_ (.A1(_0751_),
    .A2(_0686_),
    .A3(_0328_),
    .A4(_0687_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3742_ (.A1(_0634_),
    .A2(_0622_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3743_ (.A1(_0749_),
    .A2(_0750_),
    .B(_0752_),
    .C(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3744_ (.A1(_0363_),
    .A2(_0372_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3745_ (.A1(_0754_),
    .A2(_0755_),
    .B(_0700_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3746_ (.I(_0504_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3747_ (.A1(_0386_),
    .A2(_0407_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3748_ (.A1(_0758_),
    .A2(_0709_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3749_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_0465_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3751_ (.A1(_0505_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3752_ (.A1(_0498_),
    .A2(_0762_),
    .B(_0698_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3753_ (.A1(_0698_),
    .A2(_0498_),
    .A3(_0762_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3754_ (.A1(_0743_),
    .A2(_0763_),
    .A3(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3755_ (.I(_0670_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3756_ (.I(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3757_ (.A1(_0689_),
    .A2(_0697_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3758_ (.A1(_0768_),
    .A2(_0701_),
    .B(_0710_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3759_ (.A1(_0761_),
    .A2(_0769_),
    .B(_0706_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3760_ (.A1(_0698_),
    .A2(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3761_ (.I(_0662_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3762_ (.A1(_0767_),
    .A2(_0771_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3763_ (.I(_2263_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3764_ (.A1(_0763_),
    .A2(_0764_),
    .B(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3765_ (.A1(_2252_),
    .A2(_2254_),
    .A3(_0596_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3767_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3768_ (.I(_0614_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3769_ (.A1(_2306_),
    .A2(_0779_),
    .A3(_0615_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3770_ (.A1(_0529_),
    .A2(_0562_),
    .B(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3771_ (.I0(_0585_),
    .I1(_0704_),
    .S(_0564_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3772_ (.I(_0552_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3773_ (.I0(_0781_),
    .I1(_0782_),
    .S(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_0601_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3775_ (.A1(_0785_),
    .A2(_0580_),
    .B(_0549_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3776_ (.A1(_0550_),
    .A2(_0784_),
    .B(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3777_ (.A1(_0631_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3778_ (.I(_0608_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3779_ (.A1(_2159_),
    .A2(_2165_),
    .A3(_2170_),
    .A4(_2184_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3780_ (.A1(_0789_),
    .A2(_0790_),
    .A3(_2481_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3781_ (.A1(_0568_),
    .A2(_0582_),
    .B(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3782_ (.A1(_0608_),
    .A2(_0348_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3783_ (.A1(_0634_),
    .A2(_0793_),
    .B(_0641_),
    .C(_2185_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3784_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3785_ (.A1(_0766_),
    .A2(_0792_),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3786_ (.A1(_0788_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3787_ (.A1(_0778_),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3788_ (.A1(_0704_),
    .A2(_0499_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3789_ (.A1(_0705_),
    .A2(_0656_),
    .B1(_0659_),
    .B2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3790_ (.A1(_0648_),
    .A2(_2261_),
    .A3(_0649_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3791_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3792_ (.A1(_0597_),
    .A2(_0635_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3793_ (.I(_0683_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3794_ (.A1(_0629_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3795_ (.I(_0548_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3796_ (.A1(_0593_),
    .A2(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3797_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3798_ (.A1(_0625_),
    .A2(_0805_),
    .B1(_0808_),
    .B2(_0613_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3799_ (.A1(_0632_),
    .A2(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3800_ (.A1(_0496_),
    .A2(_0802_),
    .B1(_0574_),
    .B2(_0803_),
    .C(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3801_ (.A1(_0798_),
    .A2(_0800_),
    .A3(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3802_ (.A1(_0765_),
    .A2(_0773_),
    .B(_0775_),
    .C(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3803_ (.I(_0642_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3804_ (.A1(_0537_),
    .A2(_2308_),
    .A3(_2354_),
    .A4(_0512_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3805_ (.A1(_0538_),
    .A2(_0814_),
    .A3(_0815_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3806_ (.A1(_0719_),
    .A2(_0716_),
    .A3(_0718_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3807_ (.I(_0733_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3808_ (.A1(_0814_),
    .A2(_0730_),
    .A3(_0817_),
    .B(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3809_ (.I(_0648_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3810_ (.A1(_0820_),
    .A2(_0653_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3811_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3812_ (.A1(_0822_),
    .A2(_0538_),
    .A3(_0815_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3813_ (.I(_0651_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3814_ (.A1(_2309_),
    .A2(_0678_),
    .B(_0338_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3815_ (.I(_0615_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3816_ (.A1(_0614_),
    .A2(_0826_),
    .B(_0354_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3817_ (.A1(_0583_),
    .A2(_0825_),
    .A3(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3818_ (.I(_2379_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3819_ (.A1(_0621_),
    .A2(_0829_),
    .B(_0604_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3820_ (.I(_0614_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3821_ (.I(_0615_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3822_ (.A1(_0831_),
    .A2(_0832_),
    .B(_0325_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3823_ (.A1(_0554_),
    .A2(_0830_),
    .A3(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3824_ (.A1(_0828_),
    .A2(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3825_ (.A1(_2309_),
    .A2(_0678_),
    .B(_2527_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3826_ (.A1(_0779_),
    .A2(_0826_),
    .B(_2448_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_0836_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3828_ (.A1(_2386_),
    .A2(_2389_),
    .A3(_2399_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3829_ (.A1(_2400_),
    .A2(_0789_),
    .B(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3830_ (.A1(_0565_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_0601_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3832_ (.I(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3833_ (.I0(_0838_),
    .I1(_0841_),
    .S(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3834_ (.A1(_0627_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3835_ (.A1(_0627_),
    .A2(_0835_),
    .B(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3836_ (.A1(_0633_),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3837_ (.A1(_0594_),
    .A2(\mod.funct3[1] ),
    .A3(_2260_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3838_ (.A1(_0657_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3839_ (.I(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3840_ (.I(_0848_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3841_ (.A1(_0312_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3842_ (.I(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3843_ (.A1(_0534_),
    .A2(_0850_),
    .B1(_0853_),
    .B2(_0535_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3844_ (.A1(_0772_),
    .A2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3845_ (.A1(_0719_),
    .A2(_0824_),
    .B(_0847_),
    .C(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3846_ (.I(_0804_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3847_ (.A1(_0789_),
    .A2(_0829_),
    .B(_0476_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3848_ (.A1(_0831_),
    .A2(_0832_),
    .B(_0268_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3849_ (.A1(_0603_),
    .A2(_0858_),
    .A3(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3850_ (.A1(_0779_),
    .A2(_0826_),
    .B(_0556_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3851_ (.A1(_2267_),
    .A2(_0678_),
    .B(_0461_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3852_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3853_ (.A1(_0554_),
    .A2(_0861_),
    .A3(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3854_ (.A1(_0860_),
    .A2(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3855_ (.A1(_0789_),
    .A2(_0829_),
    .B(_0529_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3856_ (.A1(_0831_),
    .A2(_0832_),
    .B(_2306_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3857_ (.A1(_0555_),
    .A2(_0866_),
    .A3(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3858_ (.A1(_0621_),
    .A2(_0829_),
    .B(_2338_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3859_ (.A1(_0779_),
    .A2(_0826_),
    .B(_0495_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3860_ (.A1(_0869_),
    .A2(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3861_ (.A1(_0584_),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3862_ (.A1(_0857_),
    .A2(_0868_),
    .A3(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3863_ (.A1(_0594_),
    .A2(_0595_),
    .A3(_0596_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3864_ (.A1(_0629_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3865_ (.A1(_0857_),
    .A2(_0865_),
    .B(_0873_),
    .C(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3866_ (.I(_0683_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3867_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3868_ (.I(_0669_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3869_ (.A1(_0790_),
    .A2(_0878_),
    .A3(_0879_),
    .B(_0795_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3870_ (.A1(_0592_),
    .A2(_0877_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3871_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3872_ (.A1(_0831_),
    .A2(_0832_),
    .B(_0790_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3873_ (.A1(_0578_),
    .A2(_0866_),
    .A3(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3874_ (.A1(_0541_),
    .A2(_0878_),
    .A3(_0603_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3875_ (.A1(_0882_),
    .A2(_0884_),
    .B1(_0885_),
    .B2(_0766_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3876_ (.A1(_0880_),
    .A2(_0886_),
    .B(_0646_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3877_ (.A1(_0856_),
    .A2(_0876_),
    .A3(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3878_ (.A1(_0816_),
    .A2(_0819_),
    .B1(_0823_),
    .B2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3879_ (.I(_0367_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3880_ (.A1(_0608_),
    .A2(_0350_),
    .A3(_0348_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3881_ (.A1(_0609_),
    .A2(_0793_),
    .B(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3882_ (.A1(_0748_),
    .A2(_0750_),
    .B(_0892_),
    .C(_0753_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3883_ (.A1(_0609_),
    .A2(_0349_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3884_ (.A1(_0893_),
    .A2(_0894_),
    .B(_0328_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3885_ (.A1(_0890_),
    .A2(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3886_ (.A1(_0686_),
    .A2(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3887_ (.I(_0642_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3888_ (.A1(_0604_),
    .A2(_0692_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3889_ (.I(_0326_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3890_ (.A1(_0592_),
    .A2(_0622_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3891_ (.I(_0892_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3892_ (.A1(_0564_),
    .A2(_2403_),
    .A3(_0744_),
    .B(_2459_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3893_ (.A1(_0673_),
    .A2(_0622_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3894_ (.A1(_0683_),
    .A2(_0619_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3895_ (.A1(_0747_),
    .A2(_0903_),
    .B(_0904_),
    .C(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3896_ (.A1(_0901_),
    .A2(_0902_),
    .A3(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3897_ (.A1(_0900_),
    .A2(_0351_),
    .A3(_0907_),
    .B(_0694_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3898_ (.A1(_0899_),
    .A2(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3899_ (.A1(_0898_),
    .A2(_0909_),
    .B(_0818_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3900_ (.A1(_0743_),
    .A2(_0897_),
    .B(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3901_ (.A1(_0863_),
    .A2(_0870_),
    .B(_0842_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3902_ (.I(_0552_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3903_ (.A1(_0867_),
    .A2(_0869_),
    .B(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3904_ (.A1(_0808_),
    .A2(_0912_),
    .A3(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3905_ (.A1(_0785_),
    .A2(_0858_),
    .A3(_0861_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3906_ (.A1(_0783_),
    .A2(_0830_),
    .A3(_0859_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3907_ (.A1(_0916_),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3908_ (.I(_0793_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3909_ (.A1(_0634_),
    .A2(_0919_),
    .B(_0641_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3910_ (.I(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3911_ (.A1(_0921_),
    .A2(_0885_),
    .B1(_0805_),
    .B2(_0884_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3912_ (.A1(_0626_),
    .A2(_0919_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3913_ (.A1(_0794_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3914_ (.A1(_0637_),
    .A2(_0918_),
    .B(_0922_),
    .C(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3915_ (.A1(_0915_),
    .A2(_0925_),
    .B(_0778_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3916_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3917_ (.A1(_0737_),
    .A2(_0693_),
    .B(_0927_),
    .C(_0851_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3918_ (.A1(_0686_),
    .A2(_0651_),
    .B(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3919_ (.A1(_0599_),
    .A2(_0846_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3920_ (.A1(_2264_),
    .A2(_0897_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3921_ (.A1(_0911_),
    .A2(_0926_),
    .A3(_0930_),
    .A4(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3922_ (.I(_0408_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3923_ (.A1(_0503_),
    .A2(_0489_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3924_ (.A1(_0476_),
    .A2(_0486_),
    .A3(_0488_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3925_ (.A1(_0934_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3926_ (.A1(_0356_),
    .A2(_0373_),
    .B(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3927_ (.A1(_0933_),
    .A2(_0937_),
    .A3(_0504_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3928_ (.A1(_0760_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3929_ (.A1(_0689_),
    .A2(_0697_),
    .B(_0700_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3930_ (.A1(_0933_),
    .A2(_0934_),
    .A3(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3931_ (.A1(_0934_),
    .A2(_0940_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3932_ (.A1(_0759_),
    .A2(_0942_),
    .B(_0898_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3933_ (.A1(_0814_),
    .A2(_0939_),
    .B1(_0941_),
    .B2(_0943_),
    .C(_0772_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3934_ (.A1(_0709_),
    .A2(_0850_),
    .B1(_0853_),
    .B2(_0707_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3935_ (.I0(_0611_),
    .I1(_0624_),
    .S(_0843_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3936_ (.A1(_0592_),
    .A2(_0806_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3937_ (.A1(_0785_),
    .A2(_0618_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3938_ (.I(_0576_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3939_ (.I0(_0606_),
    .I1(_0567_),
    .S(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3940_ (.A1(_0947_),
    .A2(_0948_),
    .B1(_0950_),
    .B2(_0636_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3941_ (.A1(_0808_),
    .A2(_0946_),
    .B(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3942_ (.A1(_0583_),
    .A2(_0641_),
    .A3(_0791_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3943_ (.A1(_2186_),
    .A2(_0568_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3944_ (.I0(_0954_),
    .I1(_0781_),
    .S(_0553_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3945_ (.I0(_0386_),
    .I1(_0497_),
    .S(_2380_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3946_ (.I0(_0782_),
    .I1(_0956_),
    .S(_0783_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3947_ (.I0(_0955_),
    .I1(_0957_),
    .S(_0804_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3948_ (.I(_0593_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3949_ (.A1(_0570_),
    .A2(_0953_),
    .B1(_0958_),
    .B2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_0776_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3951_ (.A1(_0795_),
    .A2(_0960_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3952_ (.A1(_0933_),
    .A2(_0651_),
    .B1(_0952_),
    .B2(_0632_),
    .C(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3953_ (.A1(_2264_),
    .A2(_0939_),
    .B(_0945_),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3954_ (.A1(_0944_),
    .A2(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3955_ (.A1(_0759_),
    .A2(_0502_),
    .A3(_0936_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3956_ (.A1(_0754_),
    .A2(_0755_),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3957_ (.A1(_0501_),
    .A2(_0507_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3958_ (.I(_0714_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3959_ (.A1(_0967_),
    .A2(_0968_),
    .B(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3960_ (.A1(_0492_),
    .A2(_0508_),
    .A3(_0714_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3961_ (.A1(_0970_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3962_ (.A1(_0725_),
    .A2(_0726_),
    .B(_0511_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3963_ (.A1(_0969_),
    .A2(_0703_),
    .A3(_0713_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3964_ (.A1(_0973_),
    .A2(_0974_),
    .B(_0643_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3965_ (.A1(_0814_),
    .A2(_0972_),
    .B(_0975_),
    .C(_0772_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3966_ (.A1(_0629_),
    .A2(_0877_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3967_ (.I(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3968_ (.A1(_0785_),
    .A2(_0830_),
    .A3(_0833_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3969_ (.A1(_0577_),
    .A2(_0858_),
    .A3(_0859_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3970_ (.A1(_0979_),
    .A2(_0980_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3971_ (.A1(_0583_),
    .A2(_0861_),
    .A3(_0863_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3972_ (.A1(_0578_),
    .A2(_0871_),
    .B(_0982_),
    .C(_0882_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3973_ (.A1(_0825_),
    .A2(_0827_),
    .B(_0601_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3974_ (.A1(_0836_),
    .A2(_0837_),
    .B(_0576_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3975_ (.A1(_0626_),
    .A2(_0562_),
    .A3(_0840_),
    .A4(_0576_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3976_ (.A1(_0806_),
    .A2(_0984_),
    .A3(_0985_),
    .B(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3977_ (.A1(_0959_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3978_ (.A1(_0978_),
    .A2(_0981_),
    .B(_0983_),
    .C(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(_0509_),
    .A2(_0650_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3980_ (.A1(_0509_),
    .A2(_0659_),
    .B(_0990_),
    .C(_0656_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3981_ (.I(_0636_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3982_ (.A1(_0842_),
    .A2(_0866_),
    .A3(_0883_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3983_ (.A1(_0913_),
    .A2(_0867_),
    .A3(_0869_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3984_ (.A1(_0993_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3985_ (.A1(_0992_),
    .A2(_0995_),
    .B(_0880_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3986_ (.A1(_0961_),
    .A2(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3987_ (.A1(_0632_),
    .A2(_0989_),
    .B1(_0991_),
    .B2(_0510_),
    .C(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3988_ (.A1(_2264_),
    .A2(_0972_),
    .B(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3989_ (.A1(_0900_),
    .A2(_0327_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3990_ (.A1(_0351_),
    .A2(_0907_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3991_ (.A1(_1000_),
    .A2(_1001_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3992_ (.A1(_2500_),
    .A2(_2529_),
    .B(_0687_),
    .C(_0355_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3993_ (.A1(_1000_),
    .A2(_1003_),
    .A3(_0370_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3994_ (.A1(_0895_),
    .A2(_1004_),
    .B(_0643_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3995_ (.A1(_0898_),
    .A2(_1002_),
    .B(_1005_),
    .C(_0818_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3996_ (.A1(_0857_),
    .A2(_0955_),
    .B(_0593_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3997_ (.I0(_0361_),
    .I1(_0503_),
    .S(_2380_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3998_ (.I0(_0691_),
    .I1(_0366_),
    .S(_0564_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3999_ (.I0(_1008_),
    .I1(_1009_),
    .S(_0949_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4000_ (.A1(_0882_),
    .A2(_1010_),
    .B1(_0957_),
    .B2(_0878_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4001_ (.A1(_0575_),
    .A2(_0921_),
    .A3(_0885_),
    .B1(_1007_),
    .B2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4002_ (.A1(_0924_),
    .A2(_1012_),
    .B(_0646_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4003_ (.A1(_0900_),
    .A2(_0802_),
    .B(_0655_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4004_ (.A1(_0878_),
    .A2(_0948_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4005_ (.A1(_0857_),
    .A2(_0946_),
    .B(_1015_),
    .C(_0599_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4006_ (.A1(_0900_),
    .A2(_0853_),
    .B1(_1014_),
    .B2(_0694_),
    .C(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4007_ (.A1(_2263_),
    .A2(_0895_),
    .A3(_1004_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4008_ (.A1(_1013_),
    .A2(_1017_),
    .A3(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4009_ (.A1(_1006_),
    .A2(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4010_ (.A1(_0616_),
    .A2(_0744_),
    .A3(_0677_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4011_ (.A1(_2460_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4012_ (.A1(_0575_),
    .A2(_0642_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4013_ (.A1(_1022_),
    .A2(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4014_ (.A1(_0821_),
    .A2(_1022_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4015_ (.A1(_0677_),
    .A2(_0801_),
    .B(_0655_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4016_ (.A1(_0677_),
    .A2(_0852_),
    .B1(_1026_),
    .B2(_2449_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4017_ (.A1(_0598_),
    .A2(_0992_),
    .A3(_0948_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4018_ (.A1(_1025_),
    .A2(_1027_),
    .A3(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4019_ (.A1(_0631_),
    .A2(_0958_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4020_ (.A1(_0565_),
    .A2(_0609_),
    .B(_0623_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4021_ (.A1(_0554_),
    .A2(_0617_),
    .A3(_0620_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4022_ (.A1(_0578_),
    .A2(_1031_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4023_ (.A1(_0540_),
    .A2(_0919_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4024_ (.A1(_0569_),
    .A2(_0843_),
    .A3(_0791_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4025_ (.A1(_1034_),
    .A2(_1035_),
    .B(_0921_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4026_ (.A1(_0978_),
    .A2(_1010_),
    .B1(_1033_),
    .B2(_0636_),
    .C(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4027_ (.A1(_1030_),
    .A2(_1037_),
    .B(_0961_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4028_ (.A1(_0818_),
    .A2(_1024_),
    .B(_1029_),
    .C(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4029_ (.A1(_0356_),
    .A2(_0373_),
    .A3(_0936_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4030_ (.A1(_0756_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4031_ (.A1(_0700_),
    .A2(_0689_),
    .A3(_0697_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4032_ (.A1(_0723_),
    .A2(_0724_),
    .B(_0936_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4033_ (.A1(_1042_),
    .A2(_1043_),
    .B(_0766_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4034_ (.A1(_0671_),
    .A2(_1041_),
    .B(_1044_),
    .C(_0733_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4035_ (.A1(_0549_),
    .A2(_0993_),
    .A3(_0994_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4036_ (.A1(_0863_),
    .A2(_0870_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4037_ (.A1(_0913_),
    .A2(_0858_),
    .A3(_0861_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4038_ (.A1(_0949_),
    .A2(_1047_),
    .B(_1048_),
    .C(_0877_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4039_ (.A1(_0959_),
    .A2(_1046_),
    .A3(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4040_ (.A1(_0795_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4041_ (.A1(_0708_),
    .A2(_0654_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4042_ (.A1(_0708_),
    .A2(_0802_),
    .B(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4043_ (.A1(_0850_),
    .A2(_1053_),
    .B(_0935_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4044_ (.A1(_0807_),
    .A2(_0984_),
    .A3(_0985_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4045_ (.A1(_0569_),
    .A2(_0843_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4046_ (.A1(_0840_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4047_ (.A1(_0805_),
    .A2(_1057_),
    .B1(_0981_),
    .B2(_0882_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4048_ (.A1(_1055_),
    .A2(_1058_),
    .B(_0598_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4049_ (.A1(_1054_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4050_ (.A1(_0822_),
    .A2(_1041_),
    .B1(_1051_),
    .B2(_0646_),
    .C(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4051_ (.A1(_0548_),
    .A2(_0619_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4052_ (.A1(_0673_),
    .A2(_2525_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4053_ (.A1(_1062_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4054_ (.I(_0747_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4055_ (.A1(_0745_),
    .A2(_0746_),
    .B(_1065_),
    .C(_1063_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4056_ (.A1(_2526_),
    .A2(_1064_),
    .A3(_1066_),
    .A4(_0902_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4057_ (.A1(_0675_),
    .A2(_0685_),
    .B(_0687_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4058_ (.A1(_0901_),
    .A2(_0902_),
    .A3(_0906_),
    .B(_0669_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4059_ (.A1(_1003_),
    .A2(_0879_),
    .A3(_1067_),
    .B1(_1068_),
    .B2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4060_ (.A1(_0582_),
    .A2(_0862_),
    .A3(_0870_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4061_ (.A1(_1071_),
    .A2(_1048_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4062_ (.A1(_0807_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4063_ (.A1(_0602_),
    .A2(_0830_),
    .A3(_0859_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4064_ (.A1(_0553_),
    .A2(_0825_),
    .A3(_0833_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4065_ (.A1(_1074_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4066_ (.A1(_0947_),
    .A2(_0995_),
    .B1(_1076_),
    .B2(_0635_),
    .C(_0924_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4067_ (.A1(_1073_),
    .A2(_1077_),
    .B(_0776_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4068_ (.A1(_0338_),
    .A2(_0349_),
    .B1(_0891_),
    .B2(_0657_),
    .C(_0848_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4069_ (.A1(_0902_),
    .A2(_0801_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4070_ (.A1(_0875_),
    .A2(_0987_),
    .B(_1079_),
    .C(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4071_ (.A1(_2262_),
    .A2(_1003_),
    .A3(_1067_),
    .B(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4072_ (.A1(_0733_),
    .A2(_1070_),
    .B(_1078_),
    .C(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(_0681_),
    .A2(_0674_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4074_ (.A1(_2528_),
    .A2(_0749_),
    .A3(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4075_ (.A1(_1062_),
    .A2(_2500_),
    .B(_1063_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4076_ (.A1(_2262_),
    .A2(_1085_),
    .A3(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4077_ (.A1(_0549_),
    .A2(_0784_),
    .B(_0786_),
    .C(_0630_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4078_ (.I0(_1008_),
    .I1(_0956_),
    .S(_0582_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4079_ (.A1(_0577_),
    .A2(_1009_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4080_ (.A1(_0949_),
    .A2(_1031_),
    .B(_0881_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4081_ (.A1(_0792_),
    .A2(_1034_),
    .B(_0920_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4082_ (.A1(_0977_),
    .A2(_1089_),
    .B1(_1090_),
    .B2(_1091_),
    .C(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4083_ (.A1(_1088_),
    .A2(_1093_),
    .B(_0777_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4084_ (.A1(_0675_),
    .A2(_0849_),
    .B1(_0852_),
    .B2(_0904_),
    .C(_0732_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4085_ (.A1(_1084_),
    .A2(_0802_),
    .B1(_0803_),
    .B2(_0625_),
    .C(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4086_ (.A1(_1065_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4087_ (.A1(_1084_),
    .A2(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4088_ (.A1(_1084_),
    .A2(_1097_),
    .B(_0879_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4089_ (.A1(_0670_),
    .A2(_1085_),
    .A3(_1086_),
    .B1(_1098_),
    .B2(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4090_ (.A1(_1087_),
    .A2(_1094_),
    .A3(_1096_),
    .B1(_1100_),
    .B2(_0663_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4091_ (.A1(_0630_),
    .A2(_1046_),
    .A3(_1049_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4092_ (.A1(_0669_),
    .A2(_1034_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4093_ (.A1(_0602_),
    .A2(_0836_),
    .A3(_0827_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4094_ (.A1(_0621_),
    .A2(_0579_),
    .B(_2403_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4095_ (.A1(_0783_),
    .A2(_0837_),
    .A3(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4096_ (.A1(_1104_),
    .A2(_1106_),
    .B(_0881_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4097_ (.A1(_0977_),
    .A2(_1076_),
    .B(_1103_),
    .C(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4098_ (.A1(_1102_),
    .A2(_1108_),
    .B(_0777_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4099_ (.A1(_0803_),
    .A2(_1057_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4100_ (.A1(_0852_),
    .A2(_0679_),
    .B1(_1105_),
    .B2(_0850_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_0616_),
    .A2(_0841_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4102_ (.A1(_0821_),
    .A2(_0650_),
    .B(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4103_ (.A1(_0662_),
    .A2(_1111_),
    .A3(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4104_ (.A1(_1109_),
    .A2(_1110_),
    .A3(_1114_),
    .B1(_1112_),
    .B2(_0663_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4105_ (.A1(_0626_),
    .A2(_0553_),
    .A3(_0866_),
    .A4(_0883_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4106_ (.A1(_0806_),
    .A2(_0912_),
    .A3(_0914_),
    .B(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4107_ (.A1(_0836_),
    .A2(_0827_),
    .B(_0842_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4108_ (.A1(_0825_),
    .A2(_0833_),
    .B(_0913_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4109_ (.A1(_0540_),
    .A2(_0919_),
    .B1(_0791_),
    .B2(_0602_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4110_ (.A1(_0881_),
    .A2(_1118_),
    .A3(_1119_),
    .B1(_0920_),
    .B2(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4111_ (.A1(_0630_),
    .A2(_1117_),
    .B1(_0918_),
    .B2(_0977_),
    .C(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4112_ (.A1(_0777_),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4113_ (.A1(_0658_),
    .A2(_0684_),
    .B(_0851_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4114_ (.A1(_0804_),
    .A2(_0619_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4115_ (.A1(_1065_),
    .A2(_0650_),
    .B1(_1124_),
    .B2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4116_ (.A1(_0844_),
    .A2(_0803_),
    .B(_1126_),
    .C(_0662_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4117_ (.A1(_2460_),
    .A2(_2463_),
    .A3(_2499_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4118_ (.A1(_2263_),
    .A2(_0749_),
    .A3(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4119_ (.A1(_1065_),
    .A2(_0903_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4120_ (.A1(_2499_),
    .A2(_0680_),
    .B(_0879_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4121_ (.A1(_0749_),
    .A2(_0670_),
    .A3(_1128_),
    .B1(_1130_),
    .B2(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4122_ (.A1(_1123_),
    .A2(_1127_),
    .A3(_1129_),
    .B1(_1132_),
    .B2(_0663_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4123_ (.A1(_1083_),
    .A2(_1101_),
    .A3(_1115_),
    .A4(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4124_ (.A1(_1039_),
    .A2(_1045_),
    .A3(_1061_),
    .A4(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4125_ (.A1(_0976_),
    .A2(_0999_),
    .A3(_1020_),
    .A4(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4126_ (.A1(_0889_),
    .A2(_0932_),
    .A3(_0965_),
    .A4(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4127_ (.A1(_0509_),
    .A2(_0973_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4128_ (.A1(_0727_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4129_ (.A1(_0727_),
    .A2(_2353_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4130_ (.A1(_0970_),
    .A2(_1140_),
    .B(_2354_),
    .C(_0512_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4131_ (.A1(_0767_),
    .A2(_1141_),
    .B(_0734_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4132_ (.A1(_0767_),
    .A2(_1139_),
    .B(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4133_ (.A1(_0555_),
    .A2(_0572_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_0584_),
    .A2(_0587_),
    .B(_0992_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4135_ (.A1(_0627_),
    .A2(_0948_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4136_ (.A1(_0550_),
    .A2(_0946_),
    .B(_1146_),
    .C(_0631_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4137_ (.A1(_0808_),
    .A2(_0950_),
    .B1(_1144_),
    .B2(_1145_),
    .C(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4138_ (.A1(_0874_),
    .A2(_1148_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4139_ (.A1(_0575_),
    .A2(_0885_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4140_ (.A1(_0637_),
    .A2(_0955_),
    .B1(_1150_),
    .B2(_0898_),
    .C(_0880_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4141_ (.A1(_0778_),
    .A2(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(_0737_),
    .A2(_2311_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4143_ (.A1(_2312_),
    .A2(_0654_),
    .A3(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4144_ (.A1(_0727_),
    .A2(_0824_),
    .B1(_1141_),
    .B2(_0822_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4145_ (.A1(_1149_),
    .A2(_1152_),
    .A3(_1154_),
    .A4(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4146_ (.I(_0505_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4147_ (.A1(_0937_),
    .A2(_0504_),
    .B(_0933_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4148_ (.A1(_0706_),
    .A2(_0463_),
    .B1(_1157_),
    .B2(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4149_ (.A1(_0761_),
    .A2(_0505_),
    .A3(_0760_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4150_ (.A1(_1159_),
    .A2(_1160_),
    .B(_0671_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4151_ (.A1(_0465_),
    .A2(_0769_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4152_ (.A1(_0743_),
    .A2(_1162_),
    .B(_0734_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4153_ (.A1(_0790_),
    .A2(_0921_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4154_ (.A1(_0959_),
    .A2(_1117_),
    .B(_0953_),
    .C(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4155_ (.A1(_0844_),
    .A2(_0805_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4156_ (.A1(_0992_),
    .A2(_0865_),
    .B1(_0978_),
    .B2(_0835_),
    .C(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4157_ (.A1(_0463_),
    .A2(_0851_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4158_ (.A1(_0652_),
    .A2(_0706_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4159_ (.A1(_0778_),
    .A2(_1165_),
    .B1(_1167_),
    .B2(_0874_),
    .C(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4160_ (.A1(_0761_),
    .A2(_0824_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4161_ (.I(_0821_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4162_ (.A1(_1172_),
    .A2(_1159_),
    .A3(_1160_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4163_ (.A1(_1161_),
    .A2(_1163_),
    .B(_1171_),
    .C(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4164_ (.A1(_0604_),
    .A2(_0692_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4165_ (.A1(_0899_),
    .A2(_0896_),
    .B(_0751_),
    .C(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4166_ (.A1(_0890_),
    .A2(_0895_),
    .B(_0899_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4167_ (.A1(_0358_),
    .A2(_1177_),
    .B(_0690_),
    .C(_0270_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4168_ (.A1(_0767_),
    .A2(_1176_),
    .A3(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4169_ (.A1(_0899_),
    .A2(_0908_),
    .B(_0693_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4170_ (.A1(_0751_),
    .A2(_1180_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4171_ (.A1(_0743_),
    .A2(_1181_),
    .B(_0734_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4172_ (.A1(_1176_),
    .A2(_1178_),
    .B(_0822_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4173_ (.A1(_1056_),
    .A2(_0923_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4174_ (.A1(_0638_),
    .A2(_0947_),
    .B1(_1184_),
    .B2(_1164_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4175_ (.A1(_0784_),
    .A2(_0978_),
    .B1(_1089_),
    .B2(_0637_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4176_ (.A1(_1185_),
    .A2(_1186_),
    .B(_0961_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(_0690_),
    .A2(_0853_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4178_ (.A1(_0270_),
    .A2(_0656_),
    .B1(_0599_),
    .B2(_0628_),
    .C(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4179_ (.A1(_0751_),
    .A2(_0824_),
    .B(_1187_),
    .C(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4180_ (.A1(_1179_),
    .A2(_1182_),
    .B(_1183_),
    .C(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4181_ (.A1(_1143_),
    .A2(_1156_),
    .A3(_1174_),
    .A4(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4182_ (.A1(_0742_),
    .A2(_0813_),
    .A3(_1137_),
    .A4(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(_0738_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4184_ (.I(_2253_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4185_ (.A1(_0741_),
    .A2(_1194_),
    .B(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4186_ (.I(_0742_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4187_ (.A1(_2253_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4188_ (.A1(_1195_),
    .A2(_1193_),
    .B(_1198_),
    .C(_0738_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4189_ (.A1(_1197_),
    .A2(_0813_),
    .A3(_1137_),
    .A4(_1192_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4190_ (.A1(_0820_),
    .A2(_0742_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4191_ (.A1(_1195_),
    .A2(_1200_),
    .B(_1201_),
    .C(_0652_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4192_ (.A1(_0645_),
    .A2(_1199_),
    .A3(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4193_ (.I(_2246_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4194_ (.I(_0661_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4195_ (.A1(_1196_),
    .A2(_1203_),
    .B(_1204_),
    .C(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4196_ (.I(\mod.valid2 ),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4197_ (.A1(_2130_),
    .A2(_1206_),
    .B(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4198_ (.I(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4199_ (.I(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4200_ (.I0(\mod.ldr_hzd[4] ),
    .I1(\mod.ldr_hzd[5] ),
    .I2(\mod.ldr_hzd[6] ),
    .I3(\mod.ldr_hzd[7] ),
    .S0(_2164_),
    .S1(_2154_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4201_ (.A1(_2150_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4202_ (.I(_2187_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4203_ (.I0(\mod.ldr_hzd[0] ),
    .I1(\mod.ldr_hzd[1] ),
    .I2(\mod.ldr_hzd[2] ),
    .I3(\mod.ldr_hzd[3] ),
    .S0(_2164_),
    .S1(_2154_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4204_ (.A1(_2126_),
    .A2(_1213_),
    .B1(_1214_),
    .B2(_2181_),
    .C(_2247_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4205_ (.I(_0401_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4206_ (.I0(\mod.ldr_hzd[0] ),
    .I1(\mod.ldr_hzd[1] ),
    .I2(\mod.ldr_hzd[2] ),
    .I3(\mod.ldr_hzd[3] ),
    .S0(_1216_),
    .S1(_0428_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4207_ (.A1(_0422_),
    .A2(\mod.ldr_hzd[5] ),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4208_ (.A1(_1216_),
    .A2(\mod.ldr_hzd[4] ),
    .B(_2348_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4209_ (.A1(_2348_),
    .A2(_1216_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4210_ (.A1(\mod.ldr_hzd[7] ),
    .A2(_0394_),
    .B1(_1220_),
    .B2(\mod.ldr_hzd[6] ),
    .C(_2270_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4211_ (.A1(_1218_),
    .A2(_1219_),
    .B(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4212_ (.A1(_0423_),
    .A2(_1217_),
    .B(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4213_ (.A1(_1205_),
    .A2(_0639_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4214_ (.A1(_1212_),
    .A2(_1215_),
    .B1(_1223_),
    .B2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4215_ (.I(_2421_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4216_ (.I(\mod.instr_2[3] ),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4217_ (.A1(_1226_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4218_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4219_ (.I(\mod.instr_2[4] ),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4220_ (.A1(_1230_),
    .A2(\mod.instr_2[3] ),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4221_ (.I(_2372_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4222_ (.A1(\mod.instr_2[4] ),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4223_ (.A1(\mod.instr_2[4] ),
    .A2(\mod.instr_2[3] ),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4224_ (.I(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4225_ (.A1(\mod.ldr_hzd[4] ),
    .A2(_1231_),
    .B1(_1233_),
    .B2(\mod.ldr_hzd[5] ),
    .C1(\mod.ldr_hzd[7] ),
    .C2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4226_ (.A1(\mod.instr_2[5] ),
    .A2(_1229_),
    .A3(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4227_ (.A1(\mod.ldr_hzd[3] ),
    .A2(_1235_),
    .B1(_1233_),
    .B2(\mod.ldr_hzd[1] ),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4228_ (.A1(\mod.ldr_hzd[0] ),
    .A2(_1231_),
    .B1(_1228_),
    .B2(\mod.ldr_hzd[2] ),
    .C(\mod.instr_2[5] ),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4229_ (.A1(_0661_),
    .A2(_0639_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4230_ (.A1(_1238_),
    .A2(_1239_),
    .B(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4231_ (.A1(_1237_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4232_ (.A1(_1205_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4233_ (.A1(\mod.ldr_hzd[4] ),
    .A2(\mod.ldr_hzd[5] ),
    .A3(\mod.ldr_hzd[6] ),
    .A4(\mod.ldr_hzd[7] ),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4234_ (.A1(\mod.ldr_hzd[0] ),
    .A2(\mod.ldr_hzd[1] ),
    .A3(\mod.ldr_hzd[2] ),
    .A4(\mod.ldr_hzd[3] ),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4235_ (.A1(_1244_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4236_ (.A1(_1225_),
    .A2(_1243_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4237_ (.A1(_1210_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4238_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4239_ (.A1(_1204_),
    .A2(_2129_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4240_ (.I(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4241_ (.I(\mod.pc_2[7] ),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4242_ (.I(_2349_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4243_ (.I(\mod.pc_2[6] ),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4244_ (.A1(_0422_),
    .A2(_0531_),
    .B(_2277_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4245_ (.A1(_1254_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4246_ (.I(\mod.pc_2[5] ),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4247_ (.A1(_1257_),
    .A2(_0449_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4248_ (.A1(_1257_),
    .A2(_0449_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4249_ (.I(\mod.pc_2[4] ),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4250_ (.I(_0405_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4251_ (.I(_0487_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4252_ (.A1(\mod.pc_2[3] ),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4253_ (.I(\mod.pc_2[2] ),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4254_ (.I0(_0820_),
    .I1(_2464_),
    .S(_0295_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4255_ (.I0(_0658_),
    .I1(_0311_),
    .S(_0295_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4256_ (.A1(\mod.pc_2[0] ),
    .A2(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4257_ (.A1(_0531_),
    .A2(_2453_),
    .B(_0296_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4258_ (.A1(\mod.pc_2[1] ),
    .A2(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4259_ (.A1(_2444_),
    .A2(_1268_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4260_ (.A1(\mod.pc_2[2] ),
    .A2(_1265_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4261_ (.A1(_1267_),
    .A2(_1269_),
    .B(_1270_),
    .C(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4262_ (.A1(_1264_),
    .A2(_1265_),
    .B(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4263_ (.A1(\mod.pc_2[3] ),
    .A2(_1262_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4264_ (.A1(_1260_),
    .A2(_1261_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4265_ (.A1(_1263_),
    .A2(_1273_),
    .B(_1274_),
    .C(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4266_ (.A1(_1260_),
    .A2(_1261_),
    .B(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4267_ (.A1(_1259_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4268_ (.A1(_1258_),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4269_ (.A1(\mod.pc_2[6] ),
    .A2(_1255_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4270_ (.A1(_1256_),
    .A2(_1279_),
    .B(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4271_ (.A1(_1252_),
    .A2(_1253_),
    .A3(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4272_ (.I(_1250_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4273_ (.A1(_0774_),
    .A2(_1191_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4274_ (.A1(_1283_),
    .A2(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4275_ (.A1(_1251_),
    .A2(_1282_),
    .B(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4276_ (.I(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4277_ (.I(_1210_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4278_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4279_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4280_ (.I(_1289_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4281_ (.I(_1247_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(\mod.pc[7] ),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4283_ (.A1(_1291_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4284_ (.A1(\mod.pc0[7] ),
    .A2(_1249_),
    .B1(_1287_),
    .B2(_1290_),
    .C(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(_2117_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4286_ (.A1(_2472_),
    .A2(_2480_),
    .B(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(_2118_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4288_ (.A1(_2126_),
    .A2(_2128_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_1213_),
    .A2(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4290_ (.I(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4291_ (.I(_1172_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_0652_),
    .A2(_1197_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4293_ (.A1(_1302_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4294_ (.A1(_1302_),
    .A2(_1115_),
    .B1(_1304_),
    .B2(_0740_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4295_ (.A1(_2400_),
    .A2(_1266_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(_1300_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4297_ (.A1(_1301_),
    .A2(_1305_),
    .B(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_1248_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4299_ (.I(\mod.pc0[0] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4300_ (.A1(_1225_),
    .A2(_1243_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4301_ (.A1(_1244_),
    .A2(_1245_),
    .B(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4302_ (.I(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4303_ (.A1(\mod.pc[0] ),
    .A2(_1289_),
    .A3(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4304_ (.A1(_1290_),
    .A2(_1308_),
    .B1(_1309_),
    .B2(_1310_),
    .C(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4305_ (.A1(_1298_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4306_ (.A1(_2123_),
    .A2(_1295_),
    .B(_1297_),
    .C(_1316_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4307_ (.I(_2122_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4308_ (.I(_1248_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4309_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4310_ (.I(_1208_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4311_ (.I(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4312_ (.I(_0774_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4313_ (.A1(_1045_),
    .A2(_1061_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4314_ (.A1(_1322_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4315_ (.A1(_1251_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(_1301_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4317_ (.I(\mod.pc_2[8] ),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4318_ (.I(_2278_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4319_ (.A1(\mod.pc_2[7] ),
    .A2(_1253_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4320_ (.A1(_1252_),
    .A2(_1253_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4321_ (.A1(_1329_),
    .A2(_1281_),
    .B(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4322_ (.A1(_1327_),
    .A2(_1328_),
    .A3(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_1326_),
    .A2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4324_ (.A1(_1321_),
    .A2(_1325_),
    .A3(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4325_ (.A1(\mod.pc[8] ),
    .A2(_1292_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4326_ (.A1(_1291_),
    .A2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4327_ (.A1(\mod.pc0[8] ),
    .A2(_1319_),
    .B(_1334_),
    .C(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4328_ (.I(_1289_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(_1302_),
    .A2(_1039_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4330_ (.A1(_1267_),
    .A2(_1269_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4331_ (.A1(_1300_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4332_ (.A1(_1301_),
    .A2(_1339_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4333_ (.A1(_1338_),
    .A2(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_2130_),
    .A2(_1206_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4335_ (.A1(\mod.valid2 ),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4336_ (.I(_1345_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4337_ (.I(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4338_ (.I(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4339_ (.A1(\mod.pc0[1] ),
    .A2(_1313_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(_1247_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4341_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4342_ (.A1(\mod.pc[1] ),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4343_ (.A1(_1348_),
    .A2(_1349_),
    .A3(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(_1343_),
    .A2(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(_1296_),
    .A2(_0590_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4346_ (.A1(_1317_),
    .A2(_1337_),
    .B1(_1354_),
    .B2(_0001_),
    .C(_1355_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4347_ (.I(_2119_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4348_ (.A1(_1267_),
    .A2(_1269_),
    .B(_1270_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4349_ (.A1(_1264_),
    .A2(_1265_),
    .A3(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4350_ (.I(_1250_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4351_ (.A1(_1302_),
    .A2(_1133_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4353_ (.A1(_1283_),
    .A2(_1358_),
    .B(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4354_ (.I(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4355_ (.I(_1288_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(_1247_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4357_ (.A1(\mod.pc[2] ),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4358_ (.A1(_1364_),
    .A2(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4359_ (.A1(\mod.pc0[2] ),
    .A2(_1249_),
    .B1(_1363_),
    .B2(_1290_),
    .C(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4360_ (.I(_1248_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4361_ (.I(_1359_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4362_ (.A1(_0944_),
    .A2(_0964_),
    .B(_1322_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_1370_),
    .A2(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4364_ (.I(\mod.pc_2[9] ),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4365_ (.I(_0532_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4366_ (.A1(\mod.pc_2[8] ),
    .A2(_1328_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4367_ (.A1(_1375_),
    .A2(_1331_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4368_ (.A1(_1327_),
    .A2(_1328_),
    .B(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4369_ (.A1(_1373_),
    .A2(_1374_),
    .A3(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4370_ (.A1(_1326_),
    .A2(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4371_ (.A1(_1321_),
    .A2(_1372_),
    .A3(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(\mod.pc[9] ),
    .A2(_1365_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4373_ (.A1(_1364_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4374_ (.A1(\mod.pc0[9] ),
    .A2(_1369_),
    .B(_1380_),
    .C(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4375_ (.I(_2122_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4376_ (.I(_2117_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4377_ (.A1(_0342_),
    .A2(_0347_),
    .B(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4378_ (.A1(_1356_),
    .A2(_1368_),
    .B1(_1383_),
    .B2(_1384_),
    .C(_1386_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4379_ (.I(\mod.pc[3] ),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4380_ (.I(_1313_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4381_ (.A1(_1387_),
    .A2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4382_ (.A1(_2523_),
    .A2(_1262_),
    .A3(_1273_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4383_ (.A1(_1172_),
    .A2(_1101_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4384_ (.A1(_1359_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4385_ (.A1(_1283_),
    .A2(_1390_),
    .B(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4386_ (.A1(_1348_),
    .A2(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4387_ (.A1(\mod.pc0[3] ),
    .A2(_1249_),
    .B1(_1389_),
    .B2(_1348_),
    .C(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4388_ (.A1(\mod.pc[10] ),
    .A2(_1351_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4389_ (.A1(\mod.pc0[10] ),
    .A2(_1318_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4390_ (.I(_1370_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4391_ (.I(\mod.pc_2[10] ),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4392_ (.A1(_2244_),
    .A2(_0531_),
    .B(_2277_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4393_ (.A1(\mod.pc_2[9] ),
    .A2(_1374_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4394_ (.A1(_1373_),
    .A2(_1374_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4395_ (.A1(_1401_),
    .A2(_1377_),
    .B(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4396_ (.A1(_1399_),
    .A2(_1400_),
    .A3(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4397_ (.A1(_1322_),
    .A2(_1174_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_1370_),
    .A2(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4399_ (.A1(_1398_),
    .A2(_1404_),
    .B(_1406_),
    .C(_1210_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4400_ (.A1(_1338_),
    .A2(_1396_),
    .B(_1397_),
    .C(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4401_ (.I(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4402_ (.A1(_0304_),
    .A2(_0309_),
    .B(_1385_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4403_ (.A1(_1356_),
    .A2(_1395_),
    .B1(_1409_),
    .B2(_1384_),
    .C(_1410_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4404_ (.A1(_2113_),
    .A2(\mod.des.des_counter[0] ),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4405_ (.I(_1411_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4406_ (.A1(_0288_),
    .A2(_0293_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4407_ (.A1(_1263_),
    .A2(_1273_),
    .B(_1274_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4408_ (.A1(_1260_),
    .A2(_1261_),
    .A3(_1414_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_1172_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4410_ (.A1(_1416_),
    .A2(_1083_),
    .B(_1359_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4411_ (.A1(_1283_),
    .A2(_1415_),
    .B(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4412_ (.I(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(\mod.pc[4] ),
    .A2(_1365_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4414_ (.A1(_1364_),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4415_ (.A1(\mod.pc0[4] ),
    .A2(_1369_),
    .B1(_1419_),
    .B2(_1338_),
    .C(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4416_ (.I(_2116_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(_1350_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4418_ (.A1(\mod.pc[11] ),
    .A2(_1348_),
    .A3(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4419_ (.A1(_1416_),
    .A2(_0813_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4420_ (.A1(\mod.pc_2[10] ),
    .A2(_1400_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4421_ (.A1(_1401_),
    .A2(_1377_),
    .B(_1427_),
    .C(_1402_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4422_ (.A1(_1399_),
    .A2(_1400_),
    .B(_1428_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4423_ (.A1(_2238_),
    .A2(_0409_),
    .A3(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4424_ (.A1(_1370_),
    .A2(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4425_ (.A1(_1398_),
    .A2(_1426_),
    .B(_1431_),
    .C(_1346_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4426_ (.A1(\mod.pc0[11] ),
    .A2(_1318_),
    .B(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4427_ (.A1(_1425_),
    .A2(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4428_ (.A1(_1423_),
    .A2(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4429_ (.A1(_1412_),
    .A2(_1413_),
    .B1(_1422_),
    .B2(_0001_),
    .C(_1435_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4430_ (.I(_2238_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_1436_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4432_ (.I(\mod.pc_2[11] ),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(_1436_),
    .A2(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4434_ (.A1(_1439_),
    .A2(_1429_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4435_ (.A1(_1436_),
    .A2(_1438_),
    .B(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4436_ (.A1(_1437_),
    .A2(\mod.pc_2[12] ),
    .A3(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4437_ (.A1(_0976_),
    .A2(_0999_),
    .B(_1322_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_1398_),
    .A2(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4439_ (.A1(_1398_),
    .A2(_1442_),
    .B(_1444_),
    .C(_1288_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4440_ (.I(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(\mod.pc[12] ),
    .A2(_1292_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4442_ (.A1(_1291_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4443_ (.A1(\mod.pc0[12] ),
    .A2(_1249_),
    .B(_1446_),
    .C(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4444_ (.A1(_1258_),
    .A2(_1259_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4445_ (.A1(_1277_),
    .A2(_1450_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_0774_),
    .A2(_1020_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4447_ (.A1(_1300_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4448_ (.A1(_1301_),
    .A2(_1451_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4449_ (.I(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(\mod.pc[5] ),
    .A2(_1365_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4451_ (.A1(_1364_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4452_ (.A1(\mod.pc0[5] ),
    .A2(_1369_),
    .B1(_1455_),
    .B2(_1338_),
    .C(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4453_ (.A1(_2534_),
    .A2(_2540_),
    .B(_1385_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4454_ (.A1(_1317_),
    .A2(_1449_),
    .B1(_1458_),
    .B2(_1356_),
    .C(_1459_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4455_ (.I(_1416_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4456_ (.A1(_1143_),
    .A2(_1156_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4457_ (.A1(_1460_),
    .A2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4458_ (.I(\mod.pc_2[13] ),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4459_ (.I(\mod.pc_2[12] ),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4460_ (.A1(_1436_),
    .A2(_1464_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4461_ (.A1(_1437_),
    .A2(_1464_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4462_ (.A1(_1465_),
    .A2(_1441_),
    .B(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4463_ (.A1(_1437_),
    .A2(_1463_),
    .A3(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4464_ (.A1(_1326_),
    .A2(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4465_ (.A1(_1326_),
    .A2(_1462_),
    .B(_1469_),
    .C(_1288_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4466_ (.I(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4467_ (.A1(\mod.pc[13] ),
    .A2(_1292_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4468_ (.A1(_1291_),
    .A2(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4469_ (.A1(\mod.pc0[13] ),
    .A2(_1319_),
    .B(_1471_),
    .C(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4470_ (.A1(\mod.pc[6] ),
    .A2(_1351_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4471_ (.A1(\mod.pc0[6] ),
    .A2(_1309_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4472_ (.A1(_1254_),
    .A2(_1255_),
    .A3(_1279_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4473_ (.A1(_1416_),
    .A2(_0932_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4474_ (.A1(_1251_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4475_ (.A1(_1251_),
    .A2(_1477_),
    .B(_1479_),
    .C(_1321_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4476_ (.A1(_1290_),
    .A2(_1475_),
    .B(_1476_),
    .C(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4477_ (.A1(_2118_),
    .A2(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4478_ (.A1(_0480_),
    .A2(_0485_),
    .B(_1296_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4479_ (.A1(_2123_),
    .A2(_1474_),
    .B(_1482_),
    .C(_1483_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_2118_),
    .A2(_1305_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4481_ (.A1(_0392_),
    .A2(_0403_),
    .B(_1296_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4482_ (.A1(_2123_),
    .A2(_1284_),
    .B(_1484_),
    .C(_1485_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4483_ (.A1(_0442_),
    .A2(_0447_),
    .B(_1385_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4484_ (.A1(_1298_),
    .A2(_1339_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4485_ (.A1(_2123_),
    .A2(_1324_),
    .B(_1486_),
    .C(_1487_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4486_ (.A1(_1317_),
    .A2(_1371_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4487_ (.A1(_0427_),
    .A2(_0434_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4488_ (.A1(_1412_),
    .A2(_1489_),
    .B1(_1360_),
    .B2(_2120_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4489_ (.A1(_1488_),
    .A2(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4490_ (.I(_1491_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4491_ (.A1(_1412_),
    .A2(_2346_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4492_ (.A1(_2120_),
    .A2(_1391_),
    .B1(_1405_),
    .B2(_1384_),
    .C(_1492_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4493_ (.A1(_1460_),
    .A2(_1083_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4494_ (.A1(_1411_),
    .A2(_2282_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4495_ (.A1(_1298_),
    .A2(_1493_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4496_ (.A1(_1384_),
    .A2(_1426_),
    .B(_1495_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4497_ (.A1(_1412_),
    .A2(_0516_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4498_ (.A1(_1317_),
    .A2(_1443_),
    .B1(_1452_),
    .B2(_1356_),
    .C(_1496_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4499_ (.A1(_1411_),
    .A2(_2237_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4500_ (.A1(_1423_),
    .A2(_1462_),
    .B(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4501_ (.A1(_0001_),
    .A2(_1478_),
    .B(_1498_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4502_ (.A1(_2364_),
    .A2(_2371_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4503_ (.A1(_1207_),
    .A2(_1312_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4504_ (.A1(_1213_),
    .A2(_2117_),
    .A3(_1205_),
    .A4(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4505_ (.A1(_1460_),
    .A2(_0889_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4506_ (.A1(_1423_),
    .A2(_1502_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4507_ (.A1(_2120_),
    .A2(_1499_),
    .B1(_1501_),
    .B2(_1195_),
    .C(_1503_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4508_ (.A1(_1460_),
    .A2(_1197_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4509_ (.A1(_1423_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4510_ (.A1(_2412_),
    .A2(_2420_),
    .B(_1298_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4511_ (.A1(_1501_),
    .A2(_1505_),
    .A3(_1506_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4512_ (.I(net12),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4513_ (.I(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(_1509_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4516_ (.I(\mod.instr_2[5] ),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4517_ (.A1(\mod.valid_out3 ),
    .A2(\mod.ins_ldr_3 ),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4518_ (.I0(_1510_),
    .I1(\mod.rd_3[2] ),
    .S(_1511_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4519_ (.I(_1511_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4520_ (.A1(_2375_),
    .A2(_1500_),
    .B(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4521_ (.A1(_1507_),
    .A2(_1512_),
    .A3(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4522_ (.A1(\mod.rd_3[1] ),
    .A2(_1513_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4523_ (.A1(_1226_),
    .A2(_1513_),
    .B(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4524_ (.I(_1517_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4525_ (.I(_1511_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4526_ (.A1(\mod.rd_3[0] ),
    .A2(_1513_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4527_ (.A1(_1232_),
    .A2(_1519_),
    .B(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4529_ (.A1(_1515_),
    .A2(_1518_),
    .A3(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4530_ (.I(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4531_ (.I(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4532_ (.I(_1523_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(_1299_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_1527_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4535_ (.I(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4536_ (.A1(_1529_),
    .A2(_1305_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4537_ (.A1(\mod.valid_out3 ),
    .A2(\mod.ins_ldr_3 ),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_1204_),
    .A2(_2339_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4539_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4540_ (.A1(_1531_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4541_ (.I(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4542_ (.I(_2130_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4543_ (.A1(\mod.pc_2[0] ),
    .A2(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4544_ (.I(_1531_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4545_ (.I(\mod.des.des_dout[18] ),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4546_ (.A1(_1530_),
    .A2(_1535_),
    .A3(_1537_),
    .B1(_1538_),
    .B2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4547_ (.A1(_1526_),
    .A2(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4548_ (.A1(_2387_),
    .A2(_1525_),
    .B(_1541_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(_1519_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4550_ (.I(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4551_ (.I(_1527_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4552_ (.I(_1544_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4553_ (.I(_1534_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_1527_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4555_ (.A1(_1547_),
    .A2(_1339_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4556_ (.A1(_2444_),
    .A2(_1545_),
    .B(_1546_),
    .C(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4557_ (.A1(\mod.des.des_dout[19] ),
    .A2(_1543_),
    .B(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4558_ (.I(_1550_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4559_ (.I(_1524_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4560_ (.A1(\mod.registers.r1[1] ),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4561_ (.A1(_1525_),
    .A2(_1551_),
    .B(_1553_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4562_ (.I(_1524_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(_1554_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4564_ (.I(_2130_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4565_ (.A1(_1264_),
    .A2(_1536_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4566_ (.A1(_1556_),
    .A2(_1360_),
    .B(_1546_),
    .C(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4567_ (.A1(\mod.des.des_dout[20] ),
    .A2(_1543_),
    .B(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4569_ (.I(_1524_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4570_ (.A1(\mod.registers.r1[2] ),
    .A2(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4571_ (.A1(_1555_),
    .A2(_1560_),
    .B(_1562_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(_1556_),
    .A2(_1391_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4573_ (.A1(_2523_),
    .A2(_1545_),
    .B(_1546_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4574_ (.A1(\mod.des.des_dout[21] ),
    .A2(_1543_),
    .B1(_1563_),
    .B2(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4575_ (.I(_1565_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(\mod.registers.r1[3] ),
    .A2(_1561_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4577_ (.A1(_1555_),
    .A2(_1566_),
    .B(_1567_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4578_ (.A1(_1547_),
    .A2(_1493_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4579_ (.A1(_0607_),
    .A2(_1529_),
    .B(_1546_),
    .C(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4580_ (.A1(\mod.des.des_dout[22] ),
    .A2(_1543_),
    .B(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(\mod.registers.r1[4] ),
    .A2(_1561_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4583_ (.A1(_1555_),
    .A2(_1571_),
    .B(_1572_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4584_ (.I(_1519_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4585_ (.A1(\mod.des.des_dout[23] ),
    .A2(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4586_ (.I(_1533_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4587_ (.I(_1533_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(_1257_),
    .A2(_1544_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4589_ (.A1(_1547_),
    .A2(_1452_),
    .B(_1576_),
    .C(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4590_ (.A1(_1266_),
    .A2(_1575_),
    .B(_1578_),
    .C(_1538_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4591_ (.A1(_1574_),
    .A2(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4592_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4593_ (.I(_1523_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4594_ (.I0(_1581_),
    .I1(\mod.registers.r1[5] ),
    .S(_1582_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4595_ (.I(_1583_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(\mod.des.des_dout[24] ),
    .A2(_1542_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4597_ (.I(_1531_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4598_ (.I(_1527_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4599_ (.I(_1532_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_1254_),
    .A2(_1528_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4601_ (.A1(_1586_),
    .A2(_1478_),
    .B(_1587_),
    .C(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4602_ (.A1(_1213_),
    .A2(_2247_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(_1268_),
    .A2(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4604_ (.A1(_1585_),
    .A2(_1589_),
    .A3(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4605_ (.A1(_1584_),
    .A2(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4606_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4607_ (.I0(_1594_),
    .I1(\mod.registers.r1[6] ),
    .S(_1582_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4608_ (.I(_1595_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(\mod.des.des_dout[25] ),
    .A2(_1573_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4610_ (.A1(_1252_),
    .A2(_1544_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4611_ (.A1(_1586_),
    .A2(_1284_),
    .B(_1587_),
    .C(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_1531_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4613_ (.A1(_1265_),
    .A2(_1575_),
    .B(_1598_),
    .C(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_1596_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4615_ (.I(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4616_ (.I0(_1602_),
    .I1(\mod.registers.r1[7] ),
    .S(_1554_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4617_ (.I(_1603_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(\mod.des.des_dout[26] ),
    .A2(_1573_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4619_ (.I(_1533_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4620_ (.A1(_1327_),
    .A2(_1528_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4621_ (.A1(_1586_),
    .A2(_1324_),
    .B(_1587_),
    .C(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4622_ (.A1(_1262_),
    .A2(_1605_),
    .B(_1607_),
    .C(_1585_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4623_ (.A1(_1604_),
    .A2(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4624_ (.I(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4625_ (.A1(_1582_),
    .A2(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4626_ (.A1(_0466_),
    .A2(_1525_),
    .B(_1611_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(\mod.des.des_dout[27] ),
    .A2(_1573_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4628_ (.A1(_1373_),
    .A2(_1544_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4629_ (.A1(_1547_),
    .A2(_1371_),
    .B(_1576_),
    .C(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4630_ (.A1(_1261_),
    .A2(_1575_),
    .B(_1614_),
    .C(_1599_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(_1612_),
    .A2(_1615_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4633_ (.I0(_1617_),
    .I1(\mod.registers.r1[9] ),
    .S(_1554_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_1618_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(\mod.des.des_dout[28] ),
    .A2(_1542_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(_1399_),
    .A2(_1528_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4637_ (.A1(_1586_),
    .A2(_1405_),
    .B(_1587_),
    .C(_1620_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4638_ (.A1(_0449_),
    .A2(_1576_),
    .B(_1621_),
    .C(_1585_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_1619_),
    .A2(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4640_ (.I(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4641_ (.I0(_1624_),
    .I1(\mod.registers.r1[10] ),
    .S(_1554_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4642_ (.I(_1625_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4643_ (.I(_1519_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4644_ (.A1(_1438_),
    .A2(_1529_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4645_ (.A1(_1545_),
    .A2(_1426_),
    .B(_1575_),
    .C(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4646_ (.A1(_1255_),
    .A2(_1599_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4647_ (.A1(_1535_),
    .A2(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4648_ (.A1(\mod.des.des_dout[29] ),
    .A2(_1626_),
    .B1(_1628_),
    .B2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(\mod.registers.r1[11] ),
    .A2(_1561_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4651_ (.A1(_1555_),
    .A2(_1632_),
    .B(_1633_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4652_ (.A1(_1464_),
    .A2(_1529_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4653_ (.A1(_1545_),
    .A2(_1443_),
    .B(_1605_),
    .C(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4654_ (.A1(_1253_),
    .A2(_1599_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_1535_),
    .A2(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4656_ (.A1(\mod.des.des_dout[30] ),
    .A2(_1626_),
    .B1(_1635_),
    .B2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4657_ (.I(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4658_ (.A1(\mod.registers.r1[12] ),
    .A2(_1526_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4659_ (.A1(_1552_),
    .A2(_1639_),
    .B(_1640_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_1536_),
    .A2(_1462_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4661_ (.A1(_1463_),
    .A2(_1556_),
    .B(_1605_),
    .C(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_1328_),
    .A2(_1585_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4663_ (.A1(_1535_),
    .A2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4664_ (.A1(\mod.des.des_dout[31] ),
    .A2(_1626_),
    .B1(_1642_),
    .B2(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4665_ (.I(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(\mod.registers.r1[13] ),
    .A2(_1526_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4667_ (.A1(_1552_),
    .A2(_1646_),
    .B(_1647_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4668_ (.I(\mod.des.des_dout[32] ),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4669_ (.A1(_1536_),
    .A2(_1502_),
    .A3(_1576_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4670_ (.A1(_1374_),
    .A2(_1590_),
    .B(_1542_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4671_ (.A1(_1648_),
    .A2(_1626_),
    .B1(_1649_),
    .B2(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4672_ (.I(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4673_ (.A1(_1582_),
    .A2(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4674_ (.A1(_0522_),
    .A2(_1525_),
    .B(_1653_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4675_ (.A1(_1556_),
    .A2(_1504_),
    .A3(_1605_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(_1400_),
    .A2(_1590_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4677_ (.A1(_1538_),
    .A2(_1654_),
    .A3(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4678_ (.A1(\mod.des.des_dout[33] ),
    .A2(_1538_),
    .B(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(\mod.registers.r1[15] ),
    .A2(_1526_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4681_ (.A1(_1552_),
    .A2(_1658_),
    .B(_1659_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4682_ (.I(_1540_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4683_ (.A1(_1518_),
    .A2(_1521_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(_1515_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4685_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4686_ (.I0(_1660_),
    .I1(\mod.registers.r2[0] ),
    .S(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4687_ (.I(_1664_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(_1662_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_1665_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(_1665_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4691_ (.A1(\mod.registers.r2[1] ),
    .A2(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4692_ (.A1(_1551_),
    .A2(_1666_),
    .B(_1668_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4693_ (.A1(\mod.registers.r2[2] ),
    .A2(_1667_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_1560_),
    .A2(_1666_),
    .B(_1669_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4695_ (.I(_1663_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4696_ (.I(_1665_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4697_ (.A1(\mod.registers.r2[3] ),
    .A2(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4698_ (.A1(_1566_),
    .A2(_1670_),
    .B(_1672_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4699_ (.A1(\mod.registers.r2[4] ),
    .A2(_1671_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4700_ (.A1(_1571_),
    .A2(_1670_),
    .B(_1673_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4701_ (.I(_1663_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4702_ (.I(_1662_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4703_ (.A1(_1580_),
    .A2(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4704_ (.A1(_0302_),
    .A2(_1674_),
    .B(_1676_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4705_ (.A1(_1594_),
    .A2(_1675_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4706_ (.A1(_0281_),
    .A2(_1674_),
    .B(_1677_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4707_ (.I0(_1602_),
    .I1(\mod.registers.r2[7] ),
    .S(_1663_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(_1678_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_1665_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4710_ (.A1(_1609_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4711_ (.A1(_0478_),
    .A2(_1674_),
    .B(_1680_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4712_ (.A1(_1616_),
    .A2(_1679_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4713_ (.A1(_0388_),
    .A2(_1674_),
    .B(_1681_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4714_ (.A1(_1624_),
    .A2(_1679_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4715_ (.A1(_0454_),
    .A2(_1666_),
    .B(_1682_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(\mod.registers.r2[11] ),
    .A2(_1671_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4717_ (.A1(_1632_),
    .A2(_1670_),
    .B(_1683_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4718_ (.A1(\mod.registers.r2[12] ),
    .A2(_1671_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4719_ (.A1(_1639_),
    .A2(_1670_),
    .B(_1684_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4720_ (.A1(\mod.registers.r2[13] ),
    .A2(_1675_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4721_ (.A1(_1646_),
    .A2(_1667_),
    .B(_1685_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4722_ (.A1(_1652_),
    .A2(_1679_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4723_ (.A1(_0526_),
    .A2(_1666_),
    .B(_1686_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4724_ (.A1(\mod.registers.r2[15] ),
    .A2(_1675_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4725_ (.A1(_1658_),
    .A2(_1667_),
    .B(_1687_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4726_ (.A1(_1515_),
    .A2(_1517_),
    .A3(_1522_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4727_ (.I(_1688_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4728_ (.I(_1689_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4729_ (.I(_1688_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4730_ (.A1(_1540_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4731_ (.A1(_2381_),
    .A2(_1690_),
    .B(_1692_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4732_ (.I(_1689_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4733_ (.I(_1688_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(\mod.registers.r3[1] ),
    .A2(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_1551_),
    .A2(_1693_),
    .B(_1695_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(\mod.registers.r3[2] ),
    .A2(_1694_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4737_ (.A1(_1560_),
    .A2(_1693_),
    .B(_1696_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(\mod.registers.r3[3] ),
    .A2(_1694_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_1566_),
    .A2(_1693_),
    .B(_1697_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(\mod.registers.r3[4] ),
    .A2(_1694_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4741_ (.A1(_1571_),
    .A2(_1693_),
    .B(_1698_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4742_ (.I(_1689_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4743_ (.I0(_1581_),
    .I1(\mod.registers.r3[5] ),
    .S(_1699_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4744_ (.I(_1700_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4745_ (.A1(_1593_),
    .A2(_1691_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4746_ (.A1(_0279_),
    .A2(_1690_),
    .B(_1701_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4747_ (.I0(_1602_),
    .I1(\mod.registers.r3[7] ),
    .S(_1699_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4748_ (.I(_1702_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4749_ (.I0(_1610_),
    .I1(\mod.registers.r3[8] ),
    .S(_1699_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_1703_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4751_ (.I0(_1617_),
    .I1(\mod.registers.r3[9] ),
    .S(_1699_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4752_ (.I(_1704_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4753_ (.A1(_1623_),
    .A2(_1691_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4754_ (.A1(_0451_),
    .A2(_1690_),
    .B(_1705_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_1689_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4756_ (.I(_1688_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(\mod.registers.r3[11] ),
    .A2(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4758_ (.A1(_1632_),
    .A2(_1706_),
    .B(_1708_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4759_ (.A1(\mod.registers.r3[12] ),
    .A2(_1707_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4760_ (.A1(_1639_),
    .A2(_1706_),
    .B(_1709_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4761_ (.A1(\mod.registers.r3[13] ),
    .A2(_1707_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4762_ (.A1(_1646_),
    .A2(_1706_),
    .B(_1710_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4763_ (.A1(_1652_),
    .A2(_1691_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4764_ (.A1(_0519_),
    .A2(_1690_),
    .B(_1711_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4765_ (.A1(\mod.registers.r3[15] ),
    .A2(_1707_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4766_ (.A1(_1658_),
    .A2(_1706_),
    .B(_1712_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4767_ (.I(_1521_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4768_ (.I(_1512_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4769_ (.A1(net12),
    .A2(_1714_),
    .A3(_1514_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4770_ (.A1(_1518_),
    .A2(_1715_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_1713_),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4772_ (.I(_1717_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_1718_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4774_ (.I(_1717_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_1540_),
    .A2(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4776_ (.A1(_2385_),
    .A2(_1719_),
    .B(_1721_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4777_ (.I(_1718_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4778_ (.I(_1717_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(\mod.registers.r4[1] ),
    .A2(_1723_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4780_ (.A1(_1551_),
    .A2(_1722_),
    .B(_1724_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4781_ (.A1(\mod.registers.r4[2] ),
    .A2(_1723_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4782_ (.A1(_1560_),
    .A2(_1722_),
    .B(_1725_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4783_ (.A1(\mod.registers.r4[3] ),
    .A2(_1723_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4784_ (.A1(_1566_),
    .A2(_1722_),
    .B(_1726_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4785_ (.A1(\mod.registers.r4[4] ),
    .A2(_1723_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4786_ (.A1(_1571_),
    .A2(_1722_),
    .B(_1727_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4787_ (.I(_1718_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4788_ (.I0(_1581_),
    .I1(\mod.registers.r4[5] ),
    .S(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_1729_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4790_ (.A1(_1593_),
    .A2(_1720_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4791_ (.A1(_0272_),
    .A2(_1719_),
    .B(_1730_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4792_ (.I0(_1602_),
    .I1(\mod.registers.r4[7] ),
    .S(_1728_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4793_ (.I(_1731_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4794_ (.I0(_1610_),
    .I1(\mod.registers.r4[8] ),
    .S(_1728_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4795_ (.I(_1732_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4796_ (.I0(_1617_),
    .I1(\mod.registers.r4[9] ),
    .S(_1728_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4797_ (.I(_1733_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4798_ (.A1(_1623_),
    .A2(_1720_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4799_ (.A1(_0453_),
    .A2(_1719_),
    .B(_1734_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4800_ (.I(_1718_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(_1717_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4802_ (.A1(\mod.registers.r4[11] ),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4803_ (.A1(_1632_),
    .A2(_1735_),
    .B(_1737_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4804_ (.A1(\mod.registers.r4[12] ),
    .A2(_1736_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4805_ (.A1(_1639_),
    .A2(_1735_),
    .B(_1738_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(\mod.registers.r4[13] ),
    .A2(_1736_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4807_ (.A1(_1646_),
    .A2(_1735_),
    .B(_1739_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4808_ (.A1(_1651_),
    .A2(_1720_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4809_ (.A1(_0525_),
    .A2(_1719_),
    .B(_1740_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4810_ (.A1(\mod.registers.r4[15] ),
    .A2(_1736_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4811_ (.A1(_1658_),
    .A2(_1735_),
    .B(_1741_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4812_ (.A1(_1522_),
    .A2(_1716_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4813_ (.I(_1742_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4814_ (.I0(_1660_),
    .I1(\mod.registers.r5[0] ),
    .S(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4815_ (.I(_1744_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4816_ (.I(_1742_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4817_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_1745_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(\mod.registers.r5[1] ),
    .A2(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4820_ (.A1(_1550_),
    .A2(_1746_),
    .B(_1748_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4821_ (.I(_1745_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_1745_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4823_ (.A1(\mod.registers.r5[2] ),
    .A2(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4824_ (.A1(_1559_),
    .A2(_1749_),
    .B(_1751_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4825_ (.A1(\mod.registers.r5[3] ),
    .A2(_1750_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4826_ (.A1(_1565_),
    .A2(_1749_),
    .B(_1752_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(\mod.registers.r5[4] ),
    .A2(_1750_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4828_ (.A1(_1570_),
    .A2(_1749_),
    .B(_1753_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4829_ (.I(_1743_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_1742_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4831_ (.A1(_1580_),
    .A2(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4832_ (.A1(_0300_),
    .A2(_1754_),
    .B(_1756_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_1742_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4834_ (.A1(_1593_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4835_ (.A1(_0285_),
    .A2(_1754_),
    .B(_1758_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4836_ (.A1(_1601_),
    .A2(_1757_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4837_ (.A1(_2530_),
    .A2(_1754_),
    .B(_1759_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4838_ (.A1(_1609_),
    .A2(_1757_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4839_ (.A1(_0467_),
    .A2(_1754_),
    .B(_1760_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4840_ (.A1(_1616_),
    .A2(_1757_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4841_ (.A1(_0387_),
    .A2(_1746_),
    .B(_1761_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4842_ (.A1(_1623_),
    .A2(_1743_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4843_ (.A1(_0438_),
    .A2(_1746_),
    .B(_1762_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4844_ (.A1(\mod.registers.r5[11] ),
    .A2(_1750_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4845_ (.A1(_1631_),
    .A2(_1749_),
    .B(_1763_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4846_ (.A1(\mod.registers.r5[12] ),
    .A2(_1755_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4847_ (.A1(_1638_),
    .A2(_1747_),
    .B(_1764_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4848_ (.A1(\mod.registers.r5[13] ),
    .A2(_1755_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4849_ (.A1(_1645_),
    .A2(_1747_),
    .B(_1765_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4850_ (.A1(_1651_),
    .A2(_1743_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4851_ (.A1(_0527_),
    .A2(_1746_),
    .B(_1766_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4852_ (.A1(\mod.registers.r5[15] ),
    .A2(_1755_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4853_ (.A1(_1657_),
    .A2(_1747_),
    .B(_1767_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4854_ (.A1(_1661_),
    .A2(_1715_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4856_ (.I(_1769_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4857_ (.I0(_1660_),
    .I1(\mod.registers.r6[0] ),
    .S(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4858_ (.I(_1771_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4859_ (.I(_1768_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4860_ (.I(_1772_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(_1769_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4862_ (.A1(\mod.registers.r6[1] ),
    .A2(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4863_ (.A1(_1550_),
    .A2(_1773_),
    .B(_1775_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(\mod.registers.r6[2] ),
    .A2(_1774_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4865_ (.A1(_1559_),
    .A2(_1773_),
    .B(_1776_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(_1772_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_1769_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4868_ (.A1(\mod.registers.r6[3] ),
    .A2(_1778_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4869_ (.A1(_1565_),
    .A2(_1777_),
    .B(_1779_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4870_ (.A1(\mod.registers.r6[4] ),
    .A2(_1778_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4871_ (.A1(_1570_),
    .A2(_1777_),
    .B(_1780_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4872_ (.I0(_1581_),
    .I1(\mod.registers.r6[5] ),
    .S(_1770_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4873_ (.I(_1781_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4874_ (.I0(_1594_),
    .I1(\mod.registers.r6[6] ),
    .S(_1770_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4875_ (.I(_1782_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4876_ (.I0(_1601_),
    .I1(\mod.registers.r6[7] ),
    .S(_1770_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4877_ (.I(_1783_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4878_ (.I(_1769_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4879_ (.A1(_1609_),
    .A2(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4880_ (.A1(_0469_),
    .A2(_1773_),
    .B(_1785_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4881_ (.I0(_1617_),
    .I1(\mod.registers.r6[9] ),
    .S(_1772_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4882_ (.I(_1786_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4883_ (.I0(_1624_),
    .I1(\mod.registers.r6[10] ),
    .S(_1772_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_1787_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4885_ (.A1(\mod.registers.r6[11] ),
    .A2(_1778_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4886_ (.A1(_1631_),
    .A2(_1777_),
    .B(_1788_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4887_ (.A1(\mod.registers.r6[12] ),
    .A2(_1778_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4888_ (.A1(_1638_),
    .A2(_1777_),
    .B(_1789_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4889_ (.A1(\mod.registers.r6[13] ),
    .A2(_1784_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4890_ (.A1(_1645_),
    .A2(_1774_),
    .B(_1790_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4891_ (.A1(_1651_),
    .A2(_1784_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4892_ (.A1(_0520_),
    .A2(_1773_),
    .B(_1791_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4893_ (.A1(\mod.registers.r6[15] ),
    .A2(_1784_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4894_ (.A1(_1657_),
    .A2(_1774_),
    .B(_1792_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_1507_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4896_ (.I(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_1794_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4898_ (.I(_1795_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4899_ (.I(_1795_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4900_ (.I(_1795_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4901_ (.I(_1350_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4902_ (.I(_1796_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4903_ (.A1(\mod.valid0 ),
    .A2(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4904_ (.A1(_1795_),
    .A2(_1798_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4905_ (.I(_1796_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4906_ (.I(_1351_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4907_ (.I(_1508_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4908_ (.I(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4909_ (.A1(\mod.rd_3[0] ),
    .A2(_1800_),
    .B(_1802_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4910_ (.A1(_1232_),
    .A2(_1799_),
    .B(_1803_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4911_ (.A1(\mod.rd_3[1] ),
    .A2(_1800_),
    .B(_1802_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4912_ (.A1(_1226_),
    .A2(_1799_),
    .B(_1804_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4913_ (.I(_1793_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4914_ (.I(_1313_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4915_ (.A1(_1510_),
    .A2(_1805_),
    .A3(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4916_ (.I(_1424_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4917_ (.I(_1509_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4918_ (.A1(\mod.rd_3[2] ),
    .A2(_1808_),
    .B(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4919_ (.A1(_1807_),
    .A2(_1810_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4920_ (.A1(net12),
    .A2(_1312_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4921_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4922_ (.I(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4923_ (.A1(\mod.ins_ldr_3 ),
    .A2(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4924_ (.I(_1805_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4925_ (.A1(_1240_),
    .A2(_1799_),
    .B(_1814_),
    .C(_1815_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4926_ (.A1(\mod.ri_3 ),
    .A2(_1800_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4927_ (.A1(_2190_),
    .A2(_1799_),
    .B(_1816_),
    .C(_1815_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4928_ (.A1(\mod.pc[0] ),
    .A2(_1806_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4929_ (.A1(\mod.pc_1[0] ),
    .A2(_1808_),
    .B(_1802_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4930_ (.A1(_1817_),
    .A2(_1818_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(_1388_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(\mod.pc_1[1] ),
    .A2(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_1794_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4934_ (.A1(_1352_),
    .A2(_1820_),
    .B(_1821_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4935_ (.A1(\mod.pc_1[2] ),
    .A2(_1819_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4936_ (.A1(_1366_),
    .A2(_1822_),
    .B(_1821_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4937_ (.I(_1424_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4938_ (.A1(\mod.pc[3] ),
    .A2(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4939_ (.A1(\mod.pc_1[3] ),
    .A2(_1819_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4940_ (.A1(_1824_),
    .A2(_1825_),
    .B(_1821_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4941_ (.A1(\mod.pc_1[4] ),
    .A2(_1819_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4942_ (.A1(_1420_),
    .A2(_1826_),
    .B(_1821_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_1388_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4944_ (.A1(\mod.pc_1[5] ),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_1794_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4946_ (.A1(_1456_),
    .A2(_1828_),
    .B(_1829_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4947_ (.A1(\mod.pc_1[6] ),
    .A2(_1827_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4948_ (.A1(_1475_),
    .A2(_1830_),
    .B(_1829_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(\mod.pc_1[7] ),
    .A2(_1827_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4950_ (.A1(_1293_),
    .A2(_1831_),
    .B(_1829_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4951_ (.A1(\mod.pc_1[8] ),
    .A2(_1827_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4952_ (.A1(_1335_),
    .A2(_1832_),
    .B(_1829_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4953_ (.I(_1388_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4954_ (.A1(\mod.pc_1[9] ),
    .A2(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4955_ (.I(_1794_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4956_ (.A1(_1381_),
    .A2(_1834_),
    .B(_1835_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4957_ (.A1(\mod.pc_1[10] ),
    .A2(_1833_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4958_ (.A1(_1396_),
    .A2(_1836_),
    .B(_1835_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4959_ (.A1(\mod.pc[11] ),
    .A2(_1823_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4960_ (.A1(\mod.pc_1[11] ),
    .A2(_1833_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4961_ (.A1(_1837_),
    .A2(_1838_),
    .B(_1835_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4962_ (.A1(\mod.pc_1[12] ),
    .A2(_1833_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4963_ (.A1(_1447_),
    .A2(_1839_),
    .B(_1835_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4964_ (.A1(\mod.pc_1[13] ),
    .A2(_1806_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4965_ (.I(_1805_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4966_ (.A1(_1472_),
    .A2(_1840_),
    .B(_1841_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4967_ (.I(\mod.pc[0] ),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4968_ (.I(_1369_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4969_ (.I(_1318_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4970_ (.I0(_1842_),
    .I1(_1308_),
    .S(_1320_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4971_ (.A1(_1844_),
    .A2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4972_ (.I(_1805_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4973_ (.A1(_1842_),
    .A2(_1843_),
    .B(_1846_),
    .C(_1847_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4974_ (.I(\mod.pc[1] ),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4975_ (.I0(_1848_),
    .I1(_1342_),
    .S(_1320_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4976_ (.A1(_1845_),
    .A2(_1849_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4977_ (.A1(_1845_),
    .A2(_1849_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4978_ (.A1(_1850_),
    .A2(_1851_),
    .B(_1319_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4979_ (.A1(_1848_),
    .A2(_1843_),
    .B(_1852_),
    .C(_1847_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4980_ (.I(_1793_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4981_ (.I(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4982_ (.I(\mod.pc[2] ),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4983_ (.I0(_1855_),
    .I1(_1362_),
    .S(_1320_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(_1850_),
    .A2(_1856_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4985_ (.A1(_1850_),
    .A2(_1856_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4986_ (.A1(_1309_),
    .A2(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4987_ (.A1(\mod.pc[2] ),
    .A2(_1844_),
    .B1(_1857_),
    .B2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4988_ (.A1(_1854_),
    .A2(_1860_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4989_ (.I0(_1387_),
    .I1(_1393_),
    .S(_1209_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4990_ (.A1(_1845_),
    .A2(_1849_),
    .A3(_1856_),
    .A4(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4991_ (.I(_1862_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4992_ (.A1(_1347_),
    .A2(_1312_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_1864_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4995_ (.A1(\mod.pc[3] ),
    .A2(_1866_),
    .B(_1509_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4996_ (.A1(_1859_),
    .A2(_1861_),
    .B1(_1863_),
    .B2(_1865_),
    .C(_1867_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4997_ (.I(_1866_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4998_ (.I(\mod.pc[4] ),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4999_ (.I0(_1869_),
    .I1(_1418_),
    .S(_1209_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5000_ (.A1(_1863_),
    .A2(_1870_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5001_ (.A1(\mod.pc[4] ),
    .A2(_1865_),
    .B(_1802_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5002_ (.A1(_1868_),
    .A2(_1871_),
    .B(_1872_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5003_ (.I(\mod.pc[5] ),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5004_ (.A1(_1856_),
    .A2(_1861_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5005_ (.I0(_1873_),
    .I1(_1454_),
    .S(_1209_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5006_ (.A1(_1850_),
    .A2(_1874_),
    .A3(_1870_),
    .B(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5007_ (.A1(_1870_),
    .A2(_1875_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5008_ (.A1(_1863_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5009_ (.A1(_1876_),
    .A2(_1878_),
    .B(_1319_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5010_ (.A1(_1873_),
    .A2(_1843_),
    .B(_1879_),
    .C(_1847_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5011_ (.I(\mod.pc[6] ),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5012_ (.A1(_1880_),
    .A2(_1210_),
    .B(_1480_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5013_ (.A1(_1878_),
    .A2(_1881_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5014_ (.I(_1864_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(_1801_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5016_ (.A1(\mod.pc[6] ),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5017_ (.A1(_1868_),
    .A2(_1882_),
    .B(_1885_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5018_ (.A1(_1863_),
    .A2(_1877_),
    .A3(_1881_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5019_ (.I0(\mod.pc[7] ),
    .I1(_1287_),
    .S(_1321_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5020_ (.A1(_1886_),
    .A2(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5021_ (.A1(\mod.pc[7] ),
    .A2(_1866_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5022_ (.A1(_1865_),
    .A2(_1888_),
    .B(_1889_),
    .C(_1847_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5023_ (.A1(_1862_),
    .A2(_1877_),
    .A3(_1881_),
    .A4(_1887_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5025_ (.A1(\mod.pc[8] ),
    .A2(_1346_),
    .B(_1334_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5026_ (.A1(_1891_),
    .A2(_1892_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5027_ (.A1(_1891_),
    .A2(_1892_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5028_ (.A1(_1883_),
    .A2(_1893_),
    .A3(_1894_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(\mod.pc[8] ),
    .A2(_1843_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5030_ (.A1(_1895_),
    .A2(_1896_),
    .B(_1841_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5031_ (.A1(\mod.pc[9] ),
    .A2(_1346_),
    .B(_1380_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5032_ (.A1(_1892_),
    .A2(_1897_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5033_ (.A1(_1891_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5034_ (.A1(_1893_),
    .A2(_1897_),
    .B(_1899_),
    .C(_1309_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5035_ (.A1(\mod.pc[9] ),
    .A2(_1844_),
    .B(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5036_ (.A1(_1854_),
    .A2(_1901_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(\mod.pc[10] ),
    .A2(_1844_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5038_ (.I(_1345_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5039_ (.A1(\mod.pc[10] ),
    .A2(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5040_ (.A1(_1407_),
    .A2(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5041_ (.A1(_1899_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5042_ (.A1(_1865_),
    .A2(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5043_ (.A1(_1902_),
    .A2(_1907_),
    .B(_1841_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5044_ (.A1(_1891_),
    .A2(_1898_),
    .A3(_1905_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5045_ (.A1(\mod.pc[11] ),
    .A2(_1903_),
    .B(_1432_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5046_ (.A1(_1908_),
    .A2(_1909_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5047_ (.A1(\mod.pc[11] ),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5048_ (.A1(_1868_),
    .A2(_1910_),
    .B(_1911_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5049_ (.A1(\mod.pc[12] ),
    .A2(_1903_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5050_ (.A1(_1890_),
    .A2(_1898_),
    .A3(_1905_),
    .A4(_1909_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5051_ (.A1(_1445_),
    .A2(_1912_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5052_ (.A1(_1913_),
    .A2(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5053_ (.A1(_1913_),
    .A2(_1914_),
    .B(_1866_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5054_ (.A1(_1800_),
    .A2(_1912_),
    .B1(_1915_),
    .B2(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5055_ (.A1(_0003_),
    .A2(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5056_ (.I(_1918_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5057_ (.A1(\mod.pc[13] ),
    .A2(_1347_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5058_ (.A1(_1470_),
    .A2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5059_ (.A1(_1915_),
    .A2(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5060_ (.A1(\mod.pc[13] ),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5061_ (.A1(_1868_),
    .A2(_1921_),
    .B(_1922_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5062_ (.A1(\mod.valid0 ),
    .A2(_1347_),
    .A3(_1811_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5063_ (.I(_1923_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5064_ (.I(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5065_ (.A1(\mod.valid1 ),
    .A2(_1806_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5066_ (.A1(_1925_),
    .A2(_1926_),
    .B(_1841_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_1224_),
    .A2(_0649_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5068_ (.A1(net19),
    .A2(_1500_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5069_ (.A1(_1500_),
    .A2(_1927_),
    .B(_1928_),
    .C(_1853_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5070_ (.A1(\mod.valid1 ),
    .A2(_1903_),
    .A3(_1811_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5071_ (.I(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5072_ (.A1(_1507_),
    .A2(_1350_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_1931_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5074_ (.I(_1932_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5075_ (.A1(\mod.valid2 ),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5076_ (.A1(_1930_),
    .A2(_1934_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5077_ (.I(\mod.instr[0] ),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5078_ (.I(_1923_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5079_ (.I(_1936_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5080_ (.A1(\mod.des.des_dout[0] ),
    .A2(_1925_),
    .B(_1884_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5081_ (.A1(_1935_),
    .A2(_1937_),
    .B(_1938_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5082_ (.I(\mod.instr[1] ),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5083_ (.I(_1924_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5084_ (.I(_1801_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5085_ (.A1(\mod.des.des_dout[1] ),
    .A2(_1940_),
    .B(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5086_ (.A1(_1939_),
    .A2(_1937_),
    .B(_1942_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5087_ (.I(\mod.instr[2] ),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5088_ (.A1(\mod.des.des_dout[2] ),
    .A2(_1940_),
    .B(_1941_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5089_ (.A1(_1943_),
    .A2(_1937_),
    .B(_1944_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5090_ (.I(\mod.instr[3] ),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5091_ (.A1(\mod.des.des_dout[3] ),
    .A2(_1940_),
    .B(_1941_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5092_ (.A1(_1945_),
    .A2(_1937_),
    .B(_1946_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5093_ (.I(\mod.instr[4] ),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(_1936_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5095_ (.A1(\mod.des.des_dout[4] ),
    .A2(_1940_),
    .B(_1941_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5096_ (.A1(_1947_),
    .A2(_1948_),
    .B(_1949_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5097_ (.I(\mod.instr[5] ),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(_1924_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5099_ (.I(_1801_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5100_ (.A1(\mod.des.des_dout[5] ),
    .A2(_1951_),
    .B(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5101_ (.A1(_1950_),
    .A2(_1948_),
    .B(_1953_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5102_ (.I(\mod.instr[6] ),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5103_ (.A1(\mod.des.des_dout[6] ),
    .A2(_1951_),
    .B(_1952_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5104_ (.A1(_1954_),
    .A2(_1948_),
    .B(_1955_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5105_ (.I(\mod.instr[7] ),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5106_ (.A1(\mod.des.des_dout[7] ),
    .A2(_1951_),
    .B(_1952_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5107_ (.A1(_1956_),
    .A2(_1948_),
    .B(_1957_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5108_ (.I(\mod.instr[8] ),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5109_ (.I(_1936_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5110_ (.A1(\mod.des.des_dout[8] ),
    .A2(_1951_),
    .B(_1952_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5111_ (.A1(_1958_),
    .A2(_1959_),
    .B(_1960_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5112_ (.I(\mod.instr[9] ),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5113_ (.I(_1923_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5114_ (.I(_1508_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5115_ (.A1(\mod.des.des_dout[9] ),
    .A2(_1962_),
    .B(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5116_ (.A1(_1961_),
    .A2(_1959_),
    .B(_1964_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5117_ (.D(_0007_),
    .RN(_0003_),
    .CLK(net147),
    .Q(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5118_ (.D(_0008_),
    .CLK(net85),
    .Q(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5119_ (.D(_0009_),
    .CLK(net36),
    .Q(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5120_ (.D(_0010_),
    .CLK(net38),
    .Q(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5121_ (.D(_0011_),
    .CLK(net49),
    .Q(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5122_ (.D(_0012_),
    .CLK(net48),
    .Q(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5123_ (.D(_0013_),
    .CLK(net82),
    .Q(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5124_ (.D(_0014_),
    .CLK(net82),
    .Q(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5125_ (.D(_0015_),
    .CLK(net81),
    .Q(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5126_ (.D(_0016_),
    .CLK(net75),
    .Q(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5127_ (.D(_0017_),
    .CLK(net72),
    .Q(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5128_ (.D(_0018_),
    .CLK(net72),
    .Q(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5129_ (.D(_0019_),
    .CLK(net54),
    .Q(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5130_ (.D(_0020_),
    .CLK(net50),
    .Q(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5131_ (.D(_0021_),
    .CLK(net36),
    .Q(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5132_ (.D(_0022_),
    .CLK(net40),
    .Q(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5133_ (.D(_0023_),
    .CLK(net50),
    .Q(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5134_ (.D(_0024_),
    .CLK(net83),
    .Q(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5135_ (.D(_0025_),
    .CLK(net36),
    .Q(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5136_ (.D(_0026_),
    .CLK(net36),
    .Q(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5137_ (.D(_0027_),
    .CLK(net51),
    .Q(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5138_ (.D(_0028_),
    .CLK(net51),
    .Q(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5139_ (.D(_0029_),
    .CLK(net79),
    .Q(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5140_ (.D(_0030_),
    .CLK(net85),
    .Q(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5141_ (.D(_0031_),
    .CLK(net83),
    .Q(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5142_ (.D(_0032_),
    .CLK(net79),
    .Q(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5143_ (.D(_0033_),
    .CLK(net78),
    .Q(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5144_ (.D(_0034_),
    .CLK(net71),
    .Q(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5145_ (.D(_0035_),
    .CLK(net56),
    .Q(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5146_ (.D(_0036_),
    .CLK(net51),
    .Q(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5147_ (.D(_0037_),
    .CLK(net37),
    .Q(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5148_ (.D(_0038_),
    .CLK(net40),
    .Q(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5149_ (.D(_0039_),
    .CLK(net37),
    .Q(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5150_ (.D(_0040_),
    .CLK(net86),
    .Q(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5151_ (.D(_0041_),
    .CLK(net38),
    .Q(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5152_ (.D(_0042_),
    .CLK(net47),
    .Q(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5153_ (.D(_0043_),
    .CLK(net48),
    .Q(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5154_ (.D(_0044_),
    .CLK(net48),
    .Q(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5155_ (.D(_0045_),
    .CLK(net75),
    .Q(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5156_ (.D(_0046_),
    .CLK(net86),
    .Q(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5157_ (.D(_0047_),
    .CLK(net81),
    .Q(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5158_ (.D(_0048_),
    .CLK(net74),
    .Q(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5159_ (.D(_0049_),
    .CLK(net72),
    .Q(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5160_ (.D(_0050_),
    .CLK(net78),
    .Q(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5161_ (.D(_0051_),
    .CLK(net53),
    .Q(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5162_ (.D(_0052_),
    .CLK(net49),
    .Q(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5163_ (.D(_0053_),
    .CLK(net38),
    .Q(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5164_ (.D(_0054_),
    .CLK(net44),
    .Q(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5165_ (.D(_0055_),
    .CLK(net47),
    .Q(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5166_ (.D(_0056_),
    .CLK(net91),
    .Q(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5167_ (.D(_0057_),
    .CLK(net47),
    .Q(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5168_ (.D(_0058_),
    .CLK(net47),
    .Q(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5169_ (.D(_0059_),
    .CLK(net53),
    .Q(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5170_ (.D(_0060_),
    .CLK(net48),
    .Q(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5171_ (.D(_0061_),
    .CLK(net74),
    .Q(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5172_ (.D(_0062_),
    .CLK(net91),
    .Q(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5173_ (.D(_0063_),
    .CLK(net81),
    .Q(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5174_ (.D(_0064_),
    .CLK(net74),
    .Q(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5175_ (.D(_0065_),
    .CLK(net72),
    .Q(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5176_ (.D(_0066_),
    .CLK(net78),
    .Q(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5177_ (.D(_0067_),
    .CLK(net56),
    .Q(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5178_ (.D(_0068_),
    .CLK(net50),
    .Q(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5179_ (.D(_0069_),
    .CLK(net37),
    .Q(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5180_ (.D(_0070_),
    .CLK(net43),
    .Q(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5181_ (.D(_0071_),
    .CLK(net50),
    .Q(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5182_ (.D(_0072_),
    .CLK(net86),
    .Q(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5183_ (.D(_0073_),
    .CLK(net41),
    .Q(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5184_ (.D(_0074_),
    .CLK(net56),
    .Q(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5185_ (.D(_0075_),
    .CLK(net65),
    .Q(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5186_ (.D(_0076_),
    .CLK(net65),
    .Q(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5187_ (.D(_0077_),
    .CLK(net87),
    .Q(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5188_ (.D(_0078_),
    .CLK(net87),
    .Q(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5189_ (.D(_0079_),
    .CLK(net87),
    .Q(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5190_ (.D(_0080_),
    .CLK(net75),
    .Q(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5191_ (.D(_0081_),
    .CLK(net71),
    .Q(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5192_ (.D(_0082_),
    .CLK(net71),
    .Q(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5193_ (.D(_0083_),
    .CLK(net56),
    .Q(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5194_ (.D(_0084_),
    .CLK(net62),
    .Q(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5195_ (.D(_0085_),
    .CLK(net43),
    .Q(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5196_ (.D(_0086_),
    .CLK(net44),
    .Q(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5197_ (.D(_0087_),
    .CLK(net43),
    .Q(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5198_ (.D(_0088_),
    .CLK(net85),
    .Q(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5199_ (.D(_0089_),
    .CLK(net41),
    .Q(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5200_ (.D(_0090_),
    .CLK(net43),
    .Q(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5201_ (.D(_0091_),
    .CLK(net61),
    .Q(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5202_ (.D(_0092_),
    .CLK(net65),
    .Q(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5203_ (.D(_0093_),
    .CLK(net74),
    .Q(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5204_ (.D(_0094_),
    .CLK(net85),
    .Q(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5205_ (.D(_0095_),
    .CLK(net81),
    .Q(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5206_ (.D(_0096_),
    .CLK(net78),
    .Q(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5207_ (.D(_0097_),
    .CLK(net40),
    .Q(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5208_ (.D(_0098_),
    .CLK(net42),
    .Q(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5209_ (.D(_0099_),
    .CLK(net68),
    .Q(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5210_ (.D(_0100_),
    .CLK(net61),
    .Q(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5211_ (.D(_0101_),
    .CLK(net41),
    .Q(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5212_ (.D(_0102_),
    .CLK(net44),
    .Q(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5213_ (.D(_0103_),
    .CLK(net41),
    .Q(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5214_ (.D(_0000_),
    .SETN(_0004_),
    .CLK(net147),
    .Q(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5215_ (.D(_0001_),
    .SETN(_0005_),
    .CLK(net147),
    .Q(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5216_ (.D(_0002_),
    .SETN(_0006_),
    .CLK(net148),
    .Q(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5217_ (.D(_0104_),
    .CLK(net105),
    .Q(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5218_ (.D(_0105_),
    .CLK(net98),
    .Q(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5219_ (.D(_0106_),
    .CLK(net102),
    .Q(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5220_ (.D(_0107_),
    .CLK(net102),
    .Q(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5221_ (.D(_0108_),
    .CLK(net101),
    .Q(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5222_ (.D(_0109_),
    .CLK(net98),
    .Q(\mod.ri_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5223_ (.D(_0110_),
    .CLK(net105),
    .Q(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5224_ (.D(_0111_),
    .CLK(net129),
    .Q(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5225_ (.D(_0112_),
    .CLK(net121),
    .Q(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5226_ (.D(_0113_),
    .CLK(net128),
    .Q(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5227_ (.D(_0114_),
    .CLK(net129),
    .Q(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5228_ (.D(_0115_),
    .CLK(net129),
    .Q(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5229_ (.D(_0116_),
    .CLK(net128),
    .Q(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5230_ (.D(_0117_),
    .CLK(net128),
    .Q(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5231_ (.D(_0118_),
    .CLK(net128),
    .Q(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5232_ (.D(_0119_),
    .CLK(net119),
    .Q(\mod.pc_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5233_ (.D(_0120_),
    .CLK(net117),
    .Q(\mod.pc_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5234_ (.D(_0121_),
    .CLK(net107),
    .Q(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5235_ (.D(_0122_),
    .CLK(net107),
    .Q(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5236_ (.D(_0123_),
    .CLK(net105),
    .Q(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5237_ (.D(_0124_),
    .CLK(net109),
    .Q(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5238_ (.D(_0125_),
    .CLK(net111),
    .Q(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5239_ (.D(_0126_),
    .CLK(net120),
    .Q(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5240_ (.D(_0127_),
    .CLK(net110),
    .Q(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5241_ (.D(_0128_),
    .CLK(net109),
    .Q(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5242_ (.D(_0129_),
    .CLK(net110),
    .Q(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5243_ (.D(_0130_),
    .CLK(net109),
    .Q(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5244_ (.D(_0131_),
    .CLK(net109),
    .Q(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5245_ (.D(_0132_),
    .CLK(net110),
    .Q(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5246_ (.D(_0133_),
    .CLK(net120),
    .Q(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5247_ (.D(_0134_),
    .CLK(net106),
    .Q(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5248_ (.D(_0135_),
    .CLK(net106),
    .Q(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5249_ (.D(_0136_),
    .CLK(net106),
    .Q(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5250_ (.D(_0137_),
    .CLK(net112),
    .Q(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5251_ (.D(_0138_),
    .CLK(net102),
    .Q(\mod.valid1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5252_ (.D(_0139_),
    .CLK(net105),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5253_ (.D(_0140_),
    .CLK(net103),
    .Q(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5254_ (.D(_0141_),
    .CLK(net96),
    .Q(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5255_ (.D(_0142_),
    .CLK(net96),
    .Q(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5256_ (.D(_0143_),
    .CLK(net96),
    .Q(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5257_ (.D(_0144_),
    .CLK(net96),
    .Q(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5258_ (.D(_0145_),
    .CLK(net94),
    .Q(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5259_ (.D(_0146_),
    .CLK(net94),
    .Q(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5260_ (.D(_0147_),
    .CLK(net95),
    .Q(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5261_ (.D(_0148_),
    .CLK(net94),
    .Q(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5262_ (.D(_0149_),
    .CLK(net94),
    .Q(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5263_ (.D(_0150_),
    .CLK(net54),
    .Q(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5264_ (.D(_0151_),
    .CLK(net53),
    .Q(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5265_ (.D(_0152_),
    .CLK(net53),
    .Q(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5266_ (.D(_0153_),
    .CLK(net55),
    .Q(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5267_ (.D(_0154_),
    .CLK(net55),
    .Q(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5268_ (.D(_0155_),
    .CLK(net55),
    .Q(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5269_ (.D(_0156_),
    .CLK(net95),
    .Q(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5270_ (.D(_0157_),
    .CLK(net95),
    .Q(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5271_ (.D(_0158_),
    .CLK(net97),
    .Q(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5272_ (.D(_0159_),
    .CLK(net123),
    .Q(\mod.pc0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5273_ (.D(_0160_),
    .CLK(net120),
    .Q(\mod.pc0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5274_ (.D(_0161_),
    .CLK(net121),
    .Q(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5275_ (.D(_0162_),
    .CLK(net121),
    .Q(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5276_ (.D(_0163_),
    .CLK(net122),
    .Q(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5277_ (.D(_0164_),
    .CLK(net122),
    .Q(\mod.pc0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5278_ (.D(_0165_),
    .CLK(net120),
    .Q(\mod.pc0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5279_ (.D(_0166_),
    .CLK(net121),
    .Q(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5280_ (.D(_0167_),
    .CLK(net118),
    .Q(\mod.pc0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5281_ (.D(_0168_),
    .CLK(net118),
    .Q(\mod.pc0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5282_ (.D(_0169_),
    .CLK(net117),
    .Q(\mod.pc0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5283_ (.D(_0170_),
    .CLK(net108),
    .Q(\mod.pc0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5284_ (.D(_0171_),
    .CLK(net119),
    .Q(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5285_ (.D(_0172_),
    .CLK(net101),
    .Q(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5286_ (.D(_0173_),
    .CLK(net125),
    .Q(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5287_ (.D(_0174_),
    .CLK(net125),
    .Q(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5288_ (.D(_0175_),
    .CLK(net126),
    .Q(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5289_ (.D(_0176_),
    .CLK(net125),
    .Q(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5290_ (.D(_0177_),
    .CLK(net126),
    .Q(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5291_ (.D(_0178_),
    .CLK(net127),
    .Q(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5292_ (.D(_0179_),
    .CLK(net127),
    .Q(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5293_ (.D(_0180_),
    .CLK(net125),
    .Q(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5294_ (.D(_0181_),
    .CLK(net118),
    .Q(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5295_ (.D(_0182_),
    .CLK(net118),
    .Q(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5296_ (.D(_0183_),
    .CLK(net117),
    .Q(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5297_ (.D(_0184_),
    .CLK(net117),
    .Q(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5298_ (.D(_0185_),
    .CLK(net101),
    .Q(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5299_ (.D(_0186_),
    .CLK(net108),
    .Q(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5300_ (.D(_0187_),
    .CLK(net100),
    .Q(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5301_ (.D(_0188_),
    .CLK(net99),
    .Q(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5302_ (.D(_0189_),
    .CLK(net114),
    .Q(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5303_ (.D(_0190_),
    .CLK(net99),
    .Q(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5304_ (.D(_0191_),
    .CLK(net98),
    .Q(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5305_ (.D(_0192_),
    .CLK(net99),
    .Q(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5306_ (.D(_0193_),
    .CLK(net116),
    .Q(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5307_ (.D(_0194_),
    .CLK(net100),
    .Q(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5308_ (.D(_0195_),
    .CLK(net115),
    .Q(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5309_ (.D(_0196_),
    .CLK(net90),
    .Q(\mod.instr_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5310_ (.D(_0197_),
    .CLK(net90),
    .Q(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5311_ (.D(_0198_),
    .CLK(net67),
    .Q(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5312_ (.D(_0199_),
    .CLK(net67),
    .Q(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5313_ (.D(_0200_),
    .CLK(net90),
    .Q(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5314_ (.D(_0201_),
    .CLK(net90),
    .Q(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5315_ (.D(_0202_),
    .CLK(net114),
    .Q(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5316_ (.D(_0203_),
    .CLK(net114),
    .Q(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5317_ (.D(_0204_),
    .CLK(net114),
    .Q(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5318_ (.D(_0205_),
    .CLK(net101),
    .Q(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5319_ (.D(_0206_),
    .CLK(net66),
    .Q(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5320_ (.D(net310),
    .CLK(net57),
    .Q(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5321_ (.D(_0208_),
    .CLK(net97),
    .Q(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5322_ (.D(_0209_),
    .CLK(net66),
    .Q(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5323_ (.D(_0210_),
    .CLK(net65),
    .Q(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5324_ (.D(_0211_),
    .CLK(net98),
    .Q(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5325_ (.D(_0212_),
    .CLK(net55),
    .Q(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5326_ (.D(_0213_),
    .CLK(net66),
    .Q(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5327_ (.D(_0214_),
    .CLK(net147),
    .Q(\mod.des.des_dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5328_ (.D(_0215_),
    .CLK(net143),
    .Q(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5329_ (.D(_0216_),
    .CLK(net143),
    .Q(\mod.des.des_dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5330_ (.D(_0217_),
    .CLK(net148),
    .Q(\mod.des.des_dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5331_ (.D(_0218_),
    .CLK(net138),
    .Q(\mod.des.des_dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5332_ (.D(_0219_),
    .CLK(net138),
    .Q(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5333_ (.D(_0220_),
    .CLK(net138),
    .Q(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5334_ (.D(_0221_),
    .CLK(net136),
    .Q(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5335_ (.D(_0222_),
    .CLK(net138),
    .Q(\mod.des.des_dout[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5336_ (.D(_0223_),
    .CLK(net135),
    .Q(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5337_ (.D(_0224_),
    .CLK(net135),
    .Q(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5338_ (.D(_0225_),
    .CLK(net136),
    .Q(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5339_ (.D(_0226_),
    .CLK(net137),
    .Q(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5340_ (.D(_0227_),
    .CLK(net137),
    .Q(\mod.des.des_dout[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5341_ (.D(_0228_),
    .CLK(net136),
    .Q(\mod.des.des_dout[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5342_ (.D(_0229_),
    .CLK(net142),
    .Q(\mod.des.des_dout[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5343_ (.D(_0230_),
    .CLK(net83),
    .Q(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5344_ (.D(_0231_),
    .CLK(net62),
    .Q(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5345_ (.D(_0232_),
    .CLK(net51),
    .Q(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5346_ (.D(_0233_),
    .CLK(net60),
    .Q(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5347_ (.D(_0234_),
    .CLK(net60),
    .Q(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5348_ (.D(_0235_),
    .CLK(net76),
    .Q(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5349_ (.D(_0236_),
    .CLK(net83),
    .Q(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5350_ (.D(_0237_),
    .CLK(net84),
    .Q(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5351_ (.D(_0238_),
    .CLK(net76),
    .Q(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5352_ (.D(_0239_),
    .CLK(net73),
    .Q(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5353_ (.D(_0240_),
    .CLK(net71),
    .Q(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5354_ (.D(_0241_),
    .CLK(net60),
    .Q(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5355_ (.D(_0242_),
    .CLK(net60),
    .Q(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5356_ (.D(_0243_),
    .CLK(net62),
    .Q(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5357_ (.D(_0244_),
    .CLK(net40),
    .Q(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5358_ (.D(_0245_),
    .CLK(net62),
    .Q(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5359_ (.D(_0246_),
    .CLK(net139),
    .Q(\mod.des.des_dout[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5360_ (.D(_0247_),
    .CLK(net145),
    .Q(\mod.des.des_dout[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5361_ (.D(_0248_),
    .CLK(net139),
    .Q(\mod.des.des_dout[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5362_ (.D(_0249_),
    .CLK(net144),
    .Q(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5363_ (.D(_0250_),
    .CLK(net143),
    .Q(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5364_ (.D(_0251_),
    .CLK(net143),
    .Q(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5365_ (.D(_0252_),
    .CLK(net144),
    .Q(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5366_ (.D(_0253_),
    .CLK(net136),
    .Q(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5367_ (.D(_0254_),
    .CLK(net141),
    .Q(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5368_ (.D(_0255_),
    .CLK(net135),
    .Q(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5369_ (.D(_0256_),
    .CLK(net135),
    .Q(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5370_ (.D(_0257_),
    .CLK(net139),
    .Q(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5371_ (.D(_0258_),
    .CLK(net139),
    .Q(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5372_ (.D(_0259_),
    .CLK(net140),
    .Q(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5373_ (.D(_0260_),
    .CLK(net145),
    .Q(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5374_ (.D(_0261_),
    .CLK(net140),
    .Q(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5375_ (.D(_0262_),
    .CLK(net146),
    .Q(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5376_ (.D(_0263_),
    .CLK(net146),
    .Q(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_295 (.ZN(net295));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_296 (.ZN(net296));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_297 (.ZN(net297));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel _5320__310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(io_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input10 (.I(io_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(io_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(io_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(io_in[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(io_in[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input15 (.I(io_in[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(io_in[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(io_in[8]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(io_in[9]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout36 (.I(net39),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net46),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net42),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net45),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net45),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net45),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net70),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net52),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout50 (.I(net52),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net59),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net58),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout55 (.I(net57),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net58),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net69),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout60 (.I(net63),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net63),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout62 (.I(net64),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net68),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout65 (.I(net67),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net93),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net73),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout72 (.I(net77),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net77),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net77),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net80),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout78 (.I(net80),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net89),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout81 (.I(net84),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net84),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net88),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net92),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout90 (.I(net92),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net134),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net97),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout96 (.I(net97),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net104),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout99 (.I(net103),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout100 (.I(net103),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net103),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net113),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net107),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net111),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net111),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net111),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net133),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net116),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout116 (.I(net132),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout117 (.I(net119),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net124),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout120 (.I(net123),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout121 (.I(net123),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net131),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout125 (.I(net127),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net130),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net131),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net133),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout133 (.I(net134),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout134 (.I(\mod.clk ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout135 (.I(net137),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net142),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout138 (.I(net141),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout139 (.I(net141),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout142 (.I(net150),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout143 (.I(net145),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net149),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net149),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net149),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net1),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__RN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__D (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__D (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__D (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__B2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__B (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__B (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__C (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__B (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__B1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__B1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__I (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__I (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__C (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A3 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__B (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__B (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__C (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A3 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__B1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__B2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__B (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__B1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__B2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__B (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__C (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__B2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__B3 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A3 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A3 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__B (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I0 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__I (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__B (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__B1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__B2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I0 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__C (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A3 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A3 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A3 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__I (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A3 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A3 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A3 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A3 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A3 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A3 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A3 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__S1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A3 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A3 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A3 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A3 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A3 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__B2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__C (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A3 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A3 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A3 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__B (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__B (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__I (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A3 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__B (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A3 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A3 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A3 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A3 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__B (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__B2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__B (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__I (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__B (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__B2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__B (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A3 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__I (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__S (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__I (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__B (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__S (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__S (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__B1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A4 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__S (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__B (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__C (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__S (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I0 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__B1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__I (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__B1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__C (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__C (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__B2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A3 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__I0 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__B2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__I1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__B2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__C (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__B2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__B2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__B (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__B (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__B (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__B (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__B (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__B (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__B2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__B (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A3 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A3 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__I (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__C (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__C (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__C (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__C (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__B2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__B2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__B2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__C (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__B (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__B (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A3 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A3 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__C (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__B (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__B (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A4 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A4 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__B (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I0 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__B (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__C (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__C (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__B (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__B (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__B (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__B (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A3 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__C (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__B (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__I (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__B (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__C (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__C (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A3 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__B2 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__C (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__C (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__B (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__B (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__B (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I0 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I0 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__S (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__S (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__B (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__B1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A3 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A3 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__B (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__B (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__S (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__C (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__C (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__B (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__I0 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__B (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__B2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A3 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__C (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__I (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__C (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A3 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A3 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A3 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A3 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__B2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__C (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__B (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__B (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A3 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__C (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__B2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__C (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A4 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A3 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A3 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__B2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__B (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__B (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A4 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__B (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A3 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__B (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__C (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__C (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__B (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__B (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A3 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__S (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__S (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__B1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I0 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__B1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__C (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__B (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A3 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__C (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I0 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I0 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__C (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A3 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__B1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__C (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__C (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A3 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A3 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__B1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__B1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A3 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__B1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A3 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__B1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__B (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A3 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__C (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B2 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A3 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A3 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A4 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__B1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__C (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__B (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A3 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A3 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__B (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A4 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A4 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A3 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__C (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__C (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__B1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__S0 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__B2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__B (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__B2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A3 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__I (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__C (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__C (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__B (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__B (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__C (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__B1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A3 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__S (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__S (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__S (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__S (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__C (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__B2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A3 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__B (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__B (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__B2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__B2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__C (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__B2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A3 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__B1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__C (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__B2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__B2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__B2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__B2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__B2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__C (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__B2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__B1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__C (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__B1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__B2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__B1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__I (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__B1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__C (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__B2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__B (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__C (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__C (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__C (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__C (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__C (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A4 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__B (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I0 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__S (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__C (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__B (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__S (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__S (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__S (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__B (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__B2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A3 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__B (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I0 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I0 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I0 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__I0 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I0 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__S (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__S (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I0 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__I0 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__I0 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I0 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__I0 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A3 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__B (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__B (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__B (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I0 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I0 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__I0 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__I0 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__B (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I0 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I0 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__I0 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__B1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__B2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__B1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__B2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__B2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I0 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I0 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__I0 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I0 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I0 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__S (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__S (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__I (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__I (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__S (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__S (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__S (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__S (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A3 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__I (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__S (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__S (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__S (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__S (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__S (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__S (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__S (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__I (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A3 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A2 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__B (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__C (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__C (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__C (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A3 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__C (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__C (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__B (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__B (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__B (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__B (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__B (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__B2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A4 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__B2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__B (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A3 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A3 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A3 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__B1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__B1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__B1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__I (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__I (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__I (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__B1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__B (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__B (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__B (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__B (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__B (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__B (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__B (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__B (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__B (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__B (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__B (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__I (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__I (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__I (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__I (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__B1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__I (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__B1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__B1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A3 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__I (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__I (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__I (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__I (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__S (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__S (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__S (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__S (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__S (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__S (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__S (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__S (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__S (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__S (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__S (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__S (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__I (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__I (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__I (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__I (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__S (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__S (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__S (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__S (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__S (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__S (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__S (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__S (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__S (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__I (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__I (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__I (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__S (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__S (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__S (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__S (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__S (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__S (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__S (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__S (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__S (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__S (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__I (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__B2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__I (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__I (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__I (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__B (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__B (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__B (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__B1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__I (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__B (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__I (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__I (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__I (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__I (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A3 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A3 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A3 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A3 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A3 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A3 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__I (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__I (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__I (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__I (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__S1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__S1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A3 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A3 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A3 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__I (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A3 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A3 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A3 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__S0 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__S0 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A3 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__I (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A3 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A3 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A3 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__I (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A3 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A3 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A3 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__I (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A3 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__A3 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A3 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A3 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__I (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__I (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__B2 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__C (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__I (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__I (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__I (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__I (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__I (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__I (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__I (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A3 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A3 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A3 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A3 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__I (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A2 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__A2 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__I (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A2 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__C (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__B1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__B1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A3 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A3 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A3 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__A3 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__C1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__I (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__C1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__C1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__C1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__C1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__I (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__I (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__I (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__I (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A3 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A3 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A3 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A3 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__B1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__C1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__B1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__B1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__B1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__B1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A3 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A3 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A3 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A3 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__I (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__B1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__B1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__B1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__I (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__B (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__B2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__I (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__B2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__C (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A3 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A3 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__I (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__I (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__I (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__I (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A2 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__I (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__I (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__I (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__I (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__C (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__I (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__I (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__I (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__C (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__I (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__I (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__S (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__S (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__S (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__I (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__B (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__B (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__I (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A2 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__I (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__A3 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__I (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__I (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__I (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A3 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A3 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__A3 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__I (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__I1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A3 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A3 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A3 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A3 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A3 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A3 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__I (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A3 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A3 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A3 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__A3 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__B (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__I (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__B1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__B (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__I (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__C (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__B2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__I (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__C (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__B1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__C1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__B1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__B1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__B1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__I (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__I (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__B1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__B (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A3 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A3 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__C (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__B (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__B (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__B (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__B (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__B (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__B (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__B (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__I (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A3 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A3 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A3 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A3 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A3 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A3 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A3 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A3 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__I1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A3 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__I (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__B (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__I (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__I (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__I (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__S (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__S (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__I (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__B1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A3 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A3 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A3 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A3 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A3 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A3 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A3 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A3 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__B (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A3 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A3 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A3 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A3 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A3 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__I (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__C (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A3 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A3 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A3 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A3 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__I (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A3 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A3 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__I (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__A3 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A3 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__I (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__B (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__B (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__B (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__B2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__B (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__B1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__I (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__B1 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__B2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__I1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A3 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__I (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__I (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__I (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__I (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__B1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__I (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A3 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A3 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A3 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__B2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A3 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__I (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__B1 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__B (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__B (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__B1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A3 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A3 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A3 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A3 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__B2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A3 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__B (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__B1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__B1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__I1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A3 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A3 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__A3 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A3 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__B (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__I (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__I (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__A3 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A3 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A3 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A3 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A3 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A3 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__A3 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__I (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__B1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__I1 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__I1 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I1 (.I(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__I1 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I1 (.I(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__I1 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I1 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__I1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__I1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__I1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__I0 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__I0 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__I (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I0 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__I (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__I0 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A1 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__I (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__B2 (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__B2 (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__I (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__B2 (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__I (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__B2 (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__I (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__B2 (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__I (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__B2 (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__I (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B2 (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__I (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B2 (.I(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__I (.I(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__B2 (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__I (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__B2 (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__I (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__B2 (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__B2 (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B2 (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__B2 (.I(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__I (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B2 (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__B2 (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__B2 (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B2 (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A2 (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__I (.I(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A1 (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__I (.I(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__I (.I(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__B (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__I (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__I (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__I (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__I0 (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__I (.I(\mod.instr_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(\mod.instr_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I0 (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I0 (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B2 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I1 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I1 (.I(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A3 (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B2 (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I2 (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I2 (.I(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__I0 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__B2 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__I1 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A3 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__B2 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__I2 (.I(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A4 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__C1 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__I3 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A1 (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__I (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I (.I(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I0 (.I(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__I (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B2 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__I (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__B2 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A1 (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B2 (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B2 (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A1 (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__I (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A1 (.I(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__I (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__B2 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__I (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__B2 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__I (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__B2 (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__I (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__I (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A4 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A4 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A4 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A4 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__I (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__B2 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__I (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A4 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__B2 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__I (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__B2 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A4 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A4 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A4 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A4 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A4 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__I (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A4 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A4 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I1 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A4 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A4 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__I1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A4 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A4 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A4 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A4 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A4 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__I (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I1 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A4 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A4 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A4 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A4 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A4 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A4 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A4 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A4 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A4 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__B2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__I (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B2 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__B2 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A4 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__B2 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__A4 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__I (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A4 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__I (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__A4 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__B2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__I (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A4 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A4 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I1 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__A4 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A4 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__I (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A4 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__I (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A4 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__I (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A2 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__I (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A2 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A2 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__I (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__B2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__B2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__B2 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__C2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A2 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A2 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__I (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__B2 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__I1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A2 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A2 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__I (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__I (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A4 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A4 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A4 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__I (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A4 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__A4 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__B2 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A4 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A4 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A4 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A4 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__I (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A4 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A4 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I1 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A4 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A4 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A4 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I1 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A4 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__A4 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A4 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A4 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A4 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A4 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__I1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A4 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A4 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A4 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A4 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A4 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A4 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A4 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A4 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A4 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__I (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A4 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__I (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A4 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A4 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__I (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A4 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A4 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A4 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A4 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A4 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A4 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A4 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__A4 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__C2 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__C2 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A4 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__A4 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A4 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A4 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A4 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A4 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A4 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A4 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A4 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A4 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A4 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A4 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A4 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A4 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__I1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A4 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A4 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__I1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__I1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__I1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__I1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__I1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__I0 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__I1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__I1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__I1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__CLK (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__CLK (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__CLK (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__CLK (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__CLK (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__CLK (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__CLK (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__CLK (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__CLK (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__CLK (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__CLK (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__CLK (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1044 ();
 assign io_oeb[0] = net151;
 assign io_oeb[10] = net161;
 assign io_oeb[11] = net162;
 assign io_oeb[12] = net163;
 assign io_oeb[13] = net164;
 assign io_oeb[14] = net165;
 assign io_oeb[15] = net166;
 assign io_oeb[16] = net167;
 assign io_oeb[17] = net168;
 assign io_oeb[18] = net169;
 assign io_oeb[19] = net170;
 assign io_oeb[1] = net152;
 assign io_oeb[20] = net171;
 assign io_oeb[21] = net172;
 assign io_oeb[22] = net173;
 assign io_oeb[23] = net174;
 assign io_oeb[24] = net175;
 assign io_oeb[25] = net176;
 assign io_oeb[26] = net177;
 assign io_oeb[27] = net178;
 assign io_oeb[28] = net179;
 assign io_oeb[29] = net180;
 assign io_oeb[2] = net153;
 assign io_oeb[30] = net181;
 assign io_oeb[31] = net182;
 assign io_oeb[32] = net183;
 assign io_oeb[33] = net184;
 assign io_oeb[34] = net185;
 assign io_oeb[35] = net186;
 assign io_oeb[36] = net187;
 assign io_oeb[37] = net188;
 assign io_oeb[3] = net154;
 assign io_oeb[4] = net155;
 assign io_oeb[5] = net156;
 assign io_oeb[6] = net157;
 assign io_oeb[7] = net158;
 assign io_oeb[8] = net159;
 assign io_oeb[9] = net160;
 assign io_out[18] = net190;
 assign io_out[19] = net191;
 assign io_out[1] = net189;
 assign io_out[20] = net192;
 assign io_out[21] = net193;
 assign io_out[22] = net194;
 assign io_out[23] = net195;
 assign io_out[24] = net196;
 assign io_out[25] = net197;
 assign io_out[26] = net198;
 assign io_out[27] = net199;
 assign io_out[28] = net200;
 assign io_out[29] = net201;
 assign io_out[30] = net202;
 assign io_out[31] = net203;
 assign io_out[32] = net204;
 assign io_out[33] = net205;
 assign io_out[34] = net206;
 assign io_out[35] = net207;
 assign io_out[36] = net208;
 assign io_out[37] = net209;
 assign la_data_out[0] = net210;
 assign la_data_out[10] = net220;
 assign la_data_out[11] = net221;
 assign la_data_out[12] = net222;
 assign la_data_out[13] = net223;
 assign la_data_out[14] = net224;
 assign la_data_out[15] = net225;
 assign la_data_out[16] = net226;
 assign la_data_out[17] = net227;
 assign la_data_out[18] = net228;
 assign la_data_out[19] = net229;
 assign la_data_out[1] = net211;
 assign la_data_out[20] = net230;
 assign la_data_out[21] = net231;
 assign la_data_out[22] = net232;
 assign la_data_out[23] = net233;
 assign la_data_out[24] = net234;
 assign la_data_out[25] = net235;
 assign la_data_out[26] = net236;
 assign la_data_out[27] = net237;
 assign la_data_out[28] = net238;
 assign la_data_out[29] = net239;
 assign la_data_out[2] = net212;
 assign la_data_out[30] = net240;
 assign la_data_out[31] = net241;
 assign la_data_out[32] = net242;
 assign la_data_out[33] = net243;
 assign la_data_out[34] = net244;
 assign la_data_out[35] = net245;
 assign la_data_out[36] = net246;
 assign la_data_out[37] = net247;
 assign la_data_out[38] = net248;
 assign la_data_out[39] = net249;
 assign la_data_out[3] = net213;
 assign la_data_out[40] = net250;
 assign la_data_out[41] = net251;
 assign la_data_out[42] = net252;
 assign la_data_out[43] = net253;
 assign la_data_out[44] = net254;
 assign la_data_out[45] = net255;
 assign la_data_out[46] = net256;
 assign la_data_out[47] = net257;
 assign la_data_out[48] = net258;
 assign la_data_out[49] = net259;
 assign la_data_out[4] = net214;
 assign la_data_out[50] = net260;
 assign la_data_out[51] = net261;
 assign la_data_out[52] = net262;
 assign la_data_out[53] = net263;
 assign la_data_out[54] = net264;
 assign la_data_out[55] = net265;
 assign la_data_out[56] = net266;
 assign la_data_out[57] = net267;
 assign la_data_out[58] = net268;
 assign la_data_out[59] = net269;
 assign la_data_out[5] = net215;
 assign la_data_out[60] = net270;
 assign la_data_out[61] = net271;
 assign la_data_out[62] = net272;
 assign la_data_out[63] = net273;
 assign la_data_out[6] = net216;
 assign la_data_out[7] = net217;
 assign la_data_out[8] = net218;
 assign la_data_out[9] = net219;
 assign user_irq[0] = net274;
 assign user_irq[1] = net275;
 assign user_irq[2] = net276;
 assign wbs_ack_o = net277;
 assign wbs_dat_o[0] = net278;
 assign wbs_dat_o[10] = net288;
 assign wbs_dat_o[11] = net289;
 assign wbs_dat_o[12] = net290;
 assign wbs_dat_o[13] = net291;
 assign wbs_dat_o[14] = net292;
 assign wbs_dat_o[15] = net293;
 assign wbs_dat_o[16] = net294;
 assign wbs_dat_o[17] = net295;
 assign wbs_dat_o[18] = net296;
 assign wbs_dat_o[19] = net297;
 assign wbs_dat_o[1] = net279;
 assign wbs_dat_o[20] = net298;
 assign wbs_dat_o[21] = net299;
 assign wbs_dat_o[22] = net300;
 assign wbs_dat_o[23] = net301;
 assign wbs_dat_o[24] = net302;
 assign wbs_dat_o[25] = net303;
 assign wbs_dat_o[26] = net304;
 assign wbs_dat_o[27] = net305;
 assign wbs_dat_o[28] = net306;
 assign wbs_dat_o[29] = net307;
 assign wbs_dat_o[2] = net280;
 assign wbs_dat_o[30] = net308;
 assign wbs_dat_o[31] = net309;
 assign wbs_dat_o[3] = net281;
 assign wbs_dat_o[4] = net282;
 assign wbs_dat_o[5] = net283;
 assign wbs_dat_o[6] = net284;
 assign wbs_dat_o[7] = net285;
 assign wbs_dat_o[8] = net286;
 assign wbs_dat_o[9] = net287;
endmodule

