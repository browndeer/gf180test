// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire net217;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net218;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net219;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net255;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net274;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net275;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net276;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net277;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net278;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net279;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire \mod.clk ;
 wire \mod.des.des_counter[0] ;
 wire \mod.des.des_counter[1] ;
 wire \mod.des.des_counter[2] ;
 wire \mod.des.des_dout[0] ;
 wire \mod.des.des_dout[10] ;
 wire \mod.des.des_dout[11] ;
 wire \mod.des.des_dout[12] ;
 wire \mod.des.des_dout[13] ;
 wire \mod.des.des_dout[14] ;
 wire \mod.des.des_dout[15] ;
 wire \mod.des.des_dout[16] ;
 wire \mod.des.des_dout[17] ;
 wire \mod.des.des_dout[18] ;
 wire \mod.des.des_dout[19] ;
 wire \mod.des.des_dout[1] ;
 wire \mod.des.des_dout[20] ;
 wire \mod.des.des_dout[21] ;
 wire \mod.des.des_dout[22] ;
 wire \mod.des.des_dout[23] ;
 wire \mod.des.des_dout[24] ;
 wire \mod.des.des_dout[25] ;
 wire \mod.des.des_dout[26] ;
 wire \mod.des.des_dout[27] ;
 wire \mod.des.des_dout[28] ;
 wire \mod.des.des_dout[29] ;
 wire \mod.des.des_dout[2] ;
 wire \mod.des.des_dout[30] ;
 wire \mod.des.des_dout[31] ;
 wire \mod.des.des_dout[32] ;
 wire \mod.des.des_dout[33] ;
 wire \mod.des.des_dout[34] ;
 wire \mod.des.des_dout[35] ;
 wire \mod.des.des_dout[36] ;
 wire \mod.des.des_dout[3] ;
 wire \mod.des.des_dout[4] ;
 wire \mod.des.des_dout[5] ;
 wire \mod.des.des_dout[6] ;
 wire \mod.des.des_dout[7] ;
 wire \mod.des.des_dout[8] ;
 wire \mod.des.des_dout[9] ;
 wire \mod.funct3[0] ;
 wire \mod.funct3[1] ;
 wire \mod.funct3[2] ;
 wire \mod.funct7[0] ;
 wire \mod.funct7[1] ;
 wire \mod.funct7[2] ;
 wire \mod.ins_ldr_3 ;
 wire \mod.instr[0] ;
 wire \mod.instr[10] ;
 wire \mod.instr[11] ;
 wire \mod.instr[12] ;
 wire \mod.instr[13] ;
 wire \mod.instr[14] ;
 wire \mod.instr[15] ;
 wire \mod.instr[16] ;
 wire \mod.instr[17] ;
 wire \mod.instr[18] ;
 wire \mod.instr[19] ;
 wire \mod.instr[1] ;
 wire \mod.instr[20] ;
 wire \mod.instr[2] ;
 wire \mod.instr[3] ;
 wire \mod.instr[4] ;
 wire \mod.instr[5] ;
 wire \mod.instr[6] ;
 wire \mod.instr[7] ;
 wire \mod.instr[8] ;
 wire \mod.instr[9] ;
 wire \mod.instr_2[0] ;
 wire \mod.instr_2[10] ;
 wire \mod.instr_2[11] ;
 wire \mod.instr_2[12] ;
 wire \mod.instr_2[13] ;
 wire \mod.instr_2[14] ;
 wire \mod.instr_2[15] ;
 wire \mod.instr_2[16] ;
 wire \mod.instr_2[17] ;
 wire \mod.instr_2[1] ;
 wire \mod.instr_2[2] ;
 wire \mod.instr_2[3] ;
 wire \mod.instr_2[4] ;
 wire \mod.instr_2[5] ;
 wire \mod.instr_2[6] ;
 wire \mod.ldr_hzd[0] ;
 wire \mod.ldr_hzd[10] ;
 wire \mod.ldr_hzd[11] ;
 wire \mod.ldr_hzd[12] ;
 wire \mod.ldr_hzd[13] ;
 wire \mod.ldr_hzd[14] ;
 wire \mod.ldr_hzd[15] ;
 wire \mod.ldr_hzd[1] ;
 wire \mod.ldr_hzd[2] ;
 wire \mod.ldr_hzd[3] ;
 wire \mod.ldr_hzd[4] ;
 wire \mod.ldr_hzd[5] ;
 wire \mod.ldr_hzd[6] ;
 wire \mod.ldr_hzd[7] ;
 wire \mod.ldr_hzd[8] ;
 wire \mod.ldr_hzd[9] ;
 wire \mod.pc0[0] ;
 wire \mod.pc0[10] ;
 wire \mod.pc0[11] ;
 wire \mod.pc0[12] ;
 wire \mod.pc0[13] ;
 wire \mod.pc0[1] ;
 wire \mod.pc0[2] ;
 wire \mod.pc0[3] ;
 wire \mod.pc0[4] ;
 wire \mod.pc0[5] ;
 wire \mod.pc0[6] ;
 wire \mod.pc0[7] ;
 wire \mod.pc0[8] ;
 wire \mod.pc0[9] ;
 wire \mod.pc[0] ;
 wire \mod.pc[10] ;
 wire \mod.pc[11] ;
 wire \mod.pc[12] ;
 wire \mod.pc[13] ;
 wire \mod.pc[1] ;
 wire \mod.pc[2] ;
 wire \mod.pc[3] ;
 wire \mod.pc[4] ;
 wire \mod.pc[5] ;
 wire \mod.pc[6] ;
 wire \mod.pc[7] ;
 wire \mod.pc[8] ;
 wire \mod.pc[9] ;
 wire \mod.pc_1[0] ;
 wire \mod.pc_1[10] ;
 wire \mod.pc_1[11] ;
 wire \mod.pc_1[12] ;
 wire \mod.pc_1[13] ;
 wire \mod.pc_1[1] ;
 wire \mod.pc_1[2] ;
 wire \mod.pc_1[3] ;
 wire \mod.pc_1[4] ;
 wire \mod.pc_1[5] ;
 wire \mod.pc_1[6] ;
 wire \mod.pc_1[7] ;
 wire \mod.pc_1[8] ;
 wire \mod.pc_1[9] ;
 wire \mod.pc_2[0] ;
 wire \mod.pc_2[10] ;
 wire \mod.pc_2[11] ;
 wire \mod.pc_2[12] ;
 wire \mod.pc_2[13] ;
 wire \mod.pc_2[1] ;
 wire \mod.pc_2[2] ;
 wire \mod.pc_2[3] ;
 wire \mod.pc_2[4] ;
 wire \mod.pc_2[5] ;
 wire \mod.pc_2[6] ;
 wire \mod.pc_2[7] ;
 wire \mod.pc_2[8] ;
 wire \mod.pc_2[9] ;
 wire \mod.rd_3[0] ;
 wire \mod.rd_3[1] ;
 wire \mod.rd_3[2] ;
 wire \mod.rd_3[3] ;
 wire \mod.registers.r10[0] ;
 wire \mod.registers.r10[10] ;
 wire \mod.registers.r10[11] ;
 wire \mod.registers.r10[12] ;
 wire \mod.registers.r10[13] ;
 wire \mod.registers.r10[14] ;
 wire \mod.registers.r10[15] ;
 wire \mod.registers.r10[1] ;
 wire \mod.registers.r10[2] ;
 wire \mod.registers.r10[3] ;
 wire \mod.registers.r10[4] ;
 wire \mod.registers.r10[5] ;
 wire \mod.registers.r10[6] ;
 wire \mod.registers.r10[7] ;
 wire \mod.registers.r10[8] ;
 wire \mod.registers.r10[9] ;
 wire \mod.registers.r11[0] ;
 wire \mod.registers.r11[10] ;
 wire \mod.registers.r11[11] ;
 wire \mod.registers.r11[12] ;
 wire \mod.registers.r11[13] ;
 wire \mod.registers.r11[14] ;
 wire \mod.registers.r11[15] ;
 wire \mod.registers.r11[1] ;
 wire \mod.registers.r11[2] ;
 wire \mod.registers.r11[3] ;
 wire \mod.registers.r11[4] ;
 wire \mod.registers.r11[5] ;
 wire \mod.registers.r11[6] ;
 wire \mod.registers.r11[7] ;
 wire \mod.registers.r11[8] ;
 wire \mod.registers.r11[9] ;
 wire \mod.registers.r12[0] ;
 wire \mod.registers.r12[10] ;
 wire \mod.registers.r12[11] ;
 wire \mod.registers.r12[12] ;
 wire \mod.registers.r12[13] ;
 wire \mod.registers.r12[14] ;
 wire \mod.registers.r12[15] ;
 wire \mod.registers.r12[1] ;
 wire \mod.registers.r12[2] ;
 wire \mod.registers.r12[3] ;
 wire \mod.registers.r12[4] ;
 wire \mod.registers.r12[5] ;
 wire \mod.registers.r12[6] ;
 wire \mod.registers.r12[7] ;
 wire \mod.registers.r12[8] ;
 wire \mod.registers.r12[9] ;
 wire \mod.registers.r13[0] ;
 wire \mod.registers.r13[10] ;
 wire \mod.registers.r13[11] ;
 wire \mod.registers.r13[12] ;
 wire \mod.registers.r13[13] ;
 wire \mod.registers.r13[14] ;
 wire \mod.registers.r13[15] ;
 wire \mod.registers.r13[1] ;
 wire \mod.registers.r13[2] ;
 wire \mod.registers.r13[3] ;
 wire \mod.registers.r13[4] ;
 wire \mod.registers.r13[5] ;
 wire \mod.registers.r13[6] ;
 wire \mod.registers.r13[7] ;
 wire \mod.registers.r13[8] ;
 wire \mod.registers.r13[9] ;
 wire \mod.registers.r14[0] ;
 wire \mod.registers.r14[10] ;
 wire \mod.registers.r14[11] ;
 wire \mod.registers.r14[12] ;
 wire \mod.registers.r14[13] ;
 wire \mod.registers.r14[14] ;
 wire \mod.registers.r14[15] ;
 wire \mod.registers.r14[1] ;
 wire \mod.registers.r14[2] ;
 wire \mod.registers.r14[3] ;
 wire \mod.registers.r14[4] ;
 wire \mod.registers.r14[5] ;
 wire \mod.registers.r14[6] ;
 wire \mod.registers.r14[7] ;
 wire \mod.registers.r14[8] ;
 wire \mod.registers.r14[9] ;
 wire \mod.registers.r15[0] ;
 wire \mod.registers.r15[10] ;
 wire \mod.registers.r15[11] ;
 wire \mod.registers.r15[12] ;
 wire \mod.registers.r15[13] ;
 wire \mod.registers.r15[14] ;
 wire \mod.registers.r15[15] ;
 wire \mod.registers.r15[1] ;
 wire \mod.registers.r15[2] ;
 wire \mod.registers.r15[3] ;
 wire \mod.registers.r15[4] ;
 wire \mod.registers.r15[5] ;
 wire \mod.registers.r15[6] ;
 wire \mod.registers.r15[7] ;
 wire \mod.registers.r15[8] ;
 wire \mod.registers.r15[9] ;
 wire \mod.registers.r1[0] ;
 wire \mod.registers.r1[10] ;
 wire \mod.registers.r1[11] ;
 wire \mod.registers.r1[12] ;
 wire \mod.registers.r1[13] ;
 wire \mod.registers.r1[14] ;
 wire \mod.registers.r1[15] ;
 wire \mod.registers.r1[1] ;
 wire \mod.registers.r1[2] ;
 wire \mod.registers.r1[3] ;
 wire \mod.registers.r1[4] ;
 wire \mod.registers.r1[5] ;
 wire \mod.registers.r1[6] ;
 wire \mod.registers.r1[7] ;
 wire \mod.registers.r1[8] ;
 wire \mod.registers.r1[9] ;
 wire \mod.registers.r2[0] ;
 wire \mod.registers.r2[10] ;
 wire \mod.registers.r2[11] ;
 wire \mod.registers.r2[12] ;
 wire \mod.registers.r2[13] ;
 wire \mod.registers.r2[14] ;
 wire \mod.registers.r2[15] ;
 wire \mod.registers.r2[1] ;
 wire \mod.registers.r2[2] ;
 wire \mod.registers.r2[3] ;
 wire \mod.registers.r2[4] ;
 wire \mod.registers.r2[5] ;
 wire \mod.registers.r2[6] ;
 wire \mod.registers.r2[7] ;
 wire \mod.registers.r2[8] ;
 wire \mod.registers.r2[9] ;
 wire \mod.registers.r3[0] ;
 wire \mod.registers.r3[10] ;
 wire \mod.registers.r3[11] ;
 wire \mod.registers.r3[12] ;
 wire \mod.registers.r3[13] ;
 wire \mod.registers.r3[14] ;
 wire \mod.registers.r3[15] ;
 wire \mod.registers.r3[1] ;
 wire \mod.registers.r3[2] ;
 wire \mod.registers.r3[3] ;
 wire \mod.registers.r3[4] ;
 wire \mod.registers.r3[5] ;
 wire \mod.registers.r3[6] ;
 wire \mod.registers.r3[7] ;
 wire \mod.registers.r3[8] ;
 wire \mod.registers.r3[9] ;
 wire \mod.registers.r4[0] ;
 wire \mod.registers.r4[10] ;
 wire \mod.registers.r4[11] ;
 wire \mod.registers.r4[12] ;
 wire \mod.registers.r4[13] ;
 wire \mod.registers.r4[14] ;
 wire \mod.registers.r4[15] ;
 wire \mod.registers.r4[1] ;
 wire \mod.registers.r4[2] ;
 wire \mod.registers.r4[3] ;
 wire \mod.registers.r4[4] ;
 wire \mod.registers.r4[5] ;
 wire \mod.registers.r4[6] ;
 wire \mod.registers.r4[7] ;
 wire \mod.registers.r4[8] ;
 wire \mod.registers.r4[9] ;
 wire \mod.registers.r5[0] ;
 wire \mod.registers.r5[10] ;
 wire \mod.registers.r5[11] ;
 wire \mod.registers.r5[12] ;
 wire \mod.registers.r5[13] ;
 wire \mod.registers.r5[14] ;
 wire \mod.registers.r5[15] ;
 wire \mod.registers.r5[1] ;
 wire \mod.registers.r5[2] ;
 wire \mod.registers.r5[3] ;
 wire \mod.registers.r5[4] ;
 wire \mod.registers.r5[5] ;
 wire \mod.registers.r5[6] ;
 wire \mod.registers.r5[7] ;
 wire \mod.registers.r5[8] ;
 wire \mod.registers.r5[9] ;
 wire \mod.registers.r6[0] ;
 wire \mod.registers.r6[10] ;
 wire \mod.registers.r6[11] ;
 wire \mod.registers.r6[12] ;
 wire \mod.registers.r6[13] ;
 wire \mod.registers.r6[14] ;
 wire \mod.registers.r6[15] ;
 wire \mod.registers.r6[1] ;
 wire \mod.registers.r6[2] ;
 wire \mod.registers.r6[3] ;
 wire \mod.registers.r6[4] ;
 wire \mod.registers.r6[5] ;
 wire \mod.registers.r6[6] ;
 wire \mod.registers.r6[7] ;
 wire \mod.registers.r6[8] ;
 wire \mod.registers.r6[9] ;
 wire \mod.registers.r7[0] ;
 wire \mod.registers.r7[10] ;
 wire \mod.registers.r7[11] ;
 wire \mod.registers.r7[12] ;
 wire \mod.registers.r7[13] ;
 wire \mod.registers.r7[14] ;
 wire \mod.registers.r7[15] ;
 wire \mod.registers.r7[1] ;
 wire \mod.registers.r7[2] ;
 wire \mod.registers.r7[3] ;
 wire \mod.registers.r7[4] ;
 wire \mod.registers.r7[5] ;
 wire \mod.registers.r7[6] ;
 wire \mod.registers.r7[7] ;
 wire \mod.registers.r7[8] ;
 wire \mod.registers.r7[9] ;
 wire \mod.registers.r8[0] ;
 wire \mod.registers.r8[10] ;
 wire \mod.registers.r8[11] ;
 wire \mod.registers.r8[12] ;
 wire \mod.registers.r8[13] ;
 wire \mod.registers.r8[14] ;
 wire \mod.registers.r8[15] ;
 wire \mod.registers.r8[1] ;
 wire \mod.registers.r8[2] ;
 wire \mod.registers.r8[3] ;
 wire \mod.registers.r8[4] ;
 wire \mod.registers.r8[5] ;
 wire \mod.registers.r8[6] ;
 wire \mod.registers.r8[7] ;
 wire \mod.registers.r8[8] ;
 wire \mod.registers.r8[9] ;
 wire \mod.registers.r9[0] ;
 wire \mod.registers.r9[10] ;
 wire \mod.registers.r9[11] ;
 wire \mod.registers.r9[12] ;
 wire \mod.registers.r9[13] ;
 wire \mod.registers.r9[14] ;
 wire \mod.registers.r9[15] ;
 wire \mod.registers.r9[1] ;
 wire \mod.registers.r9[2] ;
 wire \mod.registers.r9[3] ;
 wire \mod.registers.r9[4] ;
 wire \mod.registers.r9[5] ;
 wire \mod.registers.r9[6] ;
 wire \mod.registers.r9[7] ;
 wire \mod.registers.r9[8] ;
 wire \mod.registers.r9[9] ;
 wire \mod.ri_3 ;
 wire \mod.valid0 ;
 wire \mod.valid1 ;
 wire \mod.valid2 ;
 wire \mod.valid_out3 ;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net343;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net344;
 wire net372;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3235_ (.I(\mod.des.des_counter[0] ),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3236_ (.I(\mod.des.des_counter[1] ),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3237_ (.I(_3093_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3238_ (.A1(_3092_),
    .A2(_3094_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3239_ (.A1(net141),
    .A2(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3240_ (.I(_3096_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3241_ (.I(\mod.des.des_counter[0] ),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3242_ (.I(_3097_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3243_ (.I(_3098_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3244_ (.A1(\mod.des.des_counter[0] ),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3245_ (.I(_3099_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3246_ (.I(_3100_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3247_ (.I(_3101_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3248_ (.A1(_3095_),
    .A2(_3102_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3249_ (.A1(\mod.des.des_counter[2] ),
    .A2(_3095_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3250_ (.I(_3103_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3251_ (.I(\mod.valid2 ),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3252_ (.I(_3104_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3253_ (.I(\mod.instr_2[1] ),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3254_ (.I(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3255_ (.I(_3107_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3256_ (.I(_3108_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3257_ (.I(\mod.instr_2[2] ),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3258_ (.I(_3110_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3259_ (.I(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3260_ (.I(\mod.instr_2[0] ),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3261_ (.I(_3113_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3262_ (.I(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3263_ (.A1(_3112_),
    .A2(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3264_ (.A1(_3109_),
    .A2(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3265_ (.I(\mod.funct3[1] ),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3266_ (.I(_3118_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3267_ (.I(\mod.funct3[2] ),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(_3120_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3269_ (.I(\mod.funct3[0] ),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3270_ (.A1(_3118_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3271_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3272_ (.A1(_3107_),
    .A2(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3273_ (.I(_3125_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3274_ (.I(_3126_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3275_ (.A1(_3116_),
    .A2(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3276_ (.I(_3128_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3277_ (.A1(_3121_),
    .A2(_3123_),
    .B(_3129_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3278_ (.I(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3279_ (.I(_3131_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3280_ (.I(\mod.instr_2[11] ),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3281_ (.I(_3133_),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3282_ (.I(\mod.instr_2[10] ),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3283_ (.I(_3135_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3284_ (.I(\mod.instr_2[12] ),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3285_ (.A1(\mod.instr_2[13] ),
    .A2(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3286_ (.A1(_3134_),
    .A2(_3136_),
    .A3(_3138_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3287_ (.I(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3288_ (.I(\mod.instr_2[13] ),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3289_ (.A1(_3141_),
    .A2(_3137_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3290_ (.A1(_3134_),
    .A2(_3136_),
    .A3(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3291_ (.I(_3143_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3292_ (.A1(\mod.registers.r13[7] ),
    .A2(_3140_),
    .B1(_3144_),
    .B2(\mod.registers.r1[7] ),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3293_ (.I(\mod.instr_2[13] ),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3294_ (.I(_3146_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3295_ (.I(_3137_),
    .Z(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3296_ (.A1(\mod.instr_2[11] ),
    .A2(\mod.instr_2[10] ),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3297_ (.A1(_3147_),
    .A2(_3148_),
    .A3(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3298_ (.A1(_3146_),
    .A2(_3148_),
    .A3(_3133_),
    .A4(_3135_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3299_ (.I(_3151_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3300_ (.A1(\mod.registers.r8[7] ),
    .A2(_3150_),
    .B1(_3152_),
    .B2(\mod.registers.r9[7] ),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3301_ (.I(\mod.instr_2[12] ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3302_ (.I(_3154_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3303_ (.A1(_3141_),
    .A2(_3155_),
    .A3(_3133_),
    .A4(_3135_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3304_ (.I(\mod.instr_2[11] ),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3305_ (.I(\mod.instr_2[10] ),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3306_ (.A1(_3146_),
    .A2(_3148_),
    .A3(_3157_),
    .A4(_3158_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3307_ (.I(_3159_),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3308_ (.A1(\mod.registers.r5[7] ),
    .A2(_3156_),
    .B1(_3160_),
    .B2(\mod.registers.r10[7] ),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3309_ (.A1(_3133_),
    .A2(_3158_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3310_ (.A1(_3146_),
    .A2(_3148_),
    .A3(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3311_ (.I(_3163_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3312_ (.A1(_3110_),
    .A2(_3113_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3313_ (.A1(\mod.instr_2[1] ),
    .A2(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3314_ (.I(_3166_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3315_ (.A1(\mod.registers.r11[7] ),
    .A2(_3164_),
    .B(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3316_ (.A1(_3145_),
    .A2(_3153_),
    .A3(_3161_),
    .A4(_3168_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3317_ (.A1(_3162_),
    .A2(_3142_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3318_ (.I(_3170_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3319_ (.A1(_3141_),
    .A2(_3154_),
    .A3(_3157_),
    .A4(_3158_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3320_ (.A1(\mod.registers.r3[7] ),
    .A2(_3171_),
    .B1(_3172_),
    .B2(\mod.registers.r6[7] ),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3321_ (.I(_3141_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3322_ (.I(_3149_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3323_ (.A1(_3174_),
    .A2(_3155_),
    .A3(_3175_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3324_ (.I(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3325_ (.I(_3157_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3326_ (.I(_3158_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3327_ (.A1(_3178_),
    .A2(_3179_),
    .A3(_3142_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3328_ (.I(_3180_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3329_ (.A1(\mod.registers.r4[7] ),
    .A2(_3177_),
    .B1(_3181_),
    .B2(\mod.registers.r2[7] ),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3330_ (.A1(_3178_),
    .A2(_3179_),
    .A3(_3138_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3331_ (.I(_3162_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3332_ (.A1(_3184_),
    .A2(_3138_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3333_ (.A1(\mod.registers.r14[7] ),
    .A2(_3183_),
    .B1(_3185_),
    .B2(\mod.registers.r15[7] ),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3334_ (.A1(_3174_),
    .A2(_3155_),
    .A3(_3184_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3335_ (.I(_3138_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3336_ (.A1(_3175_),
    .A2(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3337_ (.A1(\mod.registers.r7[7] ),
    .A2(_3187_),
    .B1(_3189_),
    .B2(\mod.registers.r12[7] ),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3338_ (.A1(_3173_),
    .A2(_3182_),
    .A3(_3186_),
    .A4(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3339_ (.A1(_3169_),
    .A2(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3340_ (.A1(\mod.pc_2[7] ),
    .A2(_3127_),
    .B(_3192_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3341_ (.I(\mod.funct7[2] ),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3342_ (.A1(_3194_),
    .A2(_3124_),
    .B(_3107_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3343_ (.I(_3195_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3344_ (.A1(_3110_),
    .A2(_3113_),
    .B(\mod.instr_2[1] ),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3345_ (.I(_3197_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3346_ (.I(_3198_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3347_ (.I(\mod.instr_2[17] ),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3348_ (.I(_3200_),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3349_ (.I(\mod.instr_2[16] ),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3350_ (.I(\mod.instr_2[15] ),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3351_ (.I(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3352_ (.I(\mod.instr_2[14] ),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3353_ (.A1(_3201_),
    .A2(_3202_),
    .A3(_3204_),
    .A4(_3205_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3354_ (.A1(_3200_),
    .A2(\mod.instr_2[16] ),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3355_ (.I(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3356_ (.A1(_3203_),
    .A2(\mod.instr_2[14] ),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3357_ (.A1(_3208_),
    .A2(_3209_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3358_ (.I(\mod.instr_2[15] ),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3359_ (.A1(_3211_),
    .A2(_3205_),
    .A3(_3207_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3360_ (.I(_3212_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3361_ (.A1(\mod.registers.r15[7] ),
    .A2(_3206_),
    .B1(_3210_),
    .B2(\mod.registers.r12[7] ),
    .C1(_3213_),
    .C2(\mod.registers.r14[7] ),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3362_ (.I(_3200_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3363_ (.I(\mod.instr_2[16] ),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3364_ (.I(_3216_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3365_ (.A1(_3215_),
    .A2(_3217_),
    .A3(_3209_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3366_ (.I(_3218_),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3367_ (.I(\mod.instr_2[14] ),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3368_ (.A1(_3203_),
    .A2(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3369_ (.A1(_3200_),
    .A2(_3202_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3370_ (.A1(_3221_),
    .A2(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3371_ (.I(_3223_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3372_ (.A1(_3211_),
    .A2(_3220_),
    .A3(_3222_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3373_ (.I(_3225_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3374_ (.A1(\mod.registers.r4[7] ),
    .A2(_3219_),
    .B1(_3224_),
    .B2(\mod.registers.r3[7] ),
    .C1(\mod.registers.r2[7] ),
    .C2(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3375_ (.I(\mod.instr_2[14] ),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3376_ (.I(_3228_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3377_ (.A1(_3204_),
    .A2(_3229_),
    .A3(_3222_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3378_ (.I(_3230_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3379_ (.I(_3203_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3380_ (.A1(_3232_),
    .A2(_3229_),
    .A3(_3207_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3381_ (.I(_3233_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3382_ (.A1(\mod.registers.r1[7] ),
    .A2(_3231_),
    .B1(_3234_),
    .B2(\mod.registers.r13[7] ),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3383_ (.A1(_3214_),
    .A2(_3227_),
    .A3(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3384_ (.I(\mod.instr_2[17] ),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3385_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3386_ (.I(\mod.instr_2[16] ),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3387_ (.A1(_0413_),
    .A2(_0414_),
    .A3(_3209_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3388_ (.I(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3389_ (.A1(_3201_),
    .A2(_3216_),
    .A3(_3211_),
    .A4(_3220_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3390_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3391_ (.A1(_0413_),
    .A2(_0414_),
    .A3(_3221_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3392_ (.I(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3393_ (.A1(\mod.registers.r8[7] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.registers.r6[7] ),
    .C1(_0420_),
    .C2(\mod.registers.r11[7] ),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3394_ (.A1(_3201_),
    .A2(_3217_),
    .A3(_3204_),
    .A4(_3228_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3395_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3396_ (.A1(_0412_),
    .A2(_3202_),
    .A3(_3204_),
    .A4(_3229_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3397_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3398_ (.A1(\mod.registers.r5[7] ),
    .A2(_0423_),
    .B1(_0425_),
    .B2(\mod.registers.r9[7] ),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3399_ (.I(_3211_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3400_ (.A1(_0412_),
    .A2(_0414_),
    .A3(_0427_),
    .A4(_3205_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3401_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3402_ (.A1(_3201_),
    .A2(_3217_),
    .A3(_3221_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3403_ (.I(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3404_ (.A1(\mod.registers.r10[7] ),
    .A2(_0429_),
    .B1(_0431_),
    .B2(\mod.registers.r7[7] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3405_ (.A1(_0421_),
    .A2(_0426_),
    .A3(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3406_ (.A1(_3199_),
    .A2(_0411_),
    .A3(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3407_ (.I(_3166_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3408_ (.I(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3409_ (.A1(_3110_),
    .A2(_3113_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3410_ (.A1(_0437_),
    .A2(_3197_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3411_ (.I(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3412_ (.I(\mod.instr_2[5] ),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3413_ (.I(_3217_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3414_ (.A1(\mod.funct3[2] ),
    .A2(_0437_),
    .B(_3124_),
    .C(\mod.instr_2[1] ),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3415_ (.I(_0442_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3416_ (.I0(_0440_),
    .I1(_0441_),
    .S(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3417_ (.I(_0438_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3418_ (.A1(\mod.funct3[2] ),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3419_ (.A1(_0439_),
    .A2(_0444_),
    .B(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3420_ (.A1(_0436_),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3421_ (.A1(_3196_),
    .A2(_0434_),
    .B(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3422_ (.I(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3423_ (.A1(_3193_),
    .A2(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3424_ (.I(\mod.pc_2[6] ),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3425_ (.I(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_3167_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3427_ (.I(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3429_ (.I(_3150_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3430_ (.A1(\mod.registers.r8[6] ),
    .A2(_0457_),
    .B1(_3152_),
    .B2(\mod.registers.r9[6] ),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3431_ (.A1(\mod.registers.r13[6] ),
    .A2(_3140_),
    .B1(_3144_),
    .B2(\mod.registers.r1[6] ),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3432_ (.I(_3156_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3433_ (.A1(\mod.registers.r5[6] ),
    .A2(_0460_),
    .B1(_3160_),
    .B2(\mod.registers.r10[6] ),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3434_ (.A1(\mod.registers.r11[6] ),
    .A2(_3164_),
    .B(_3167_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3435_ (.A1(_0458_),
    .A2(_0459_),
    .A3(_0461_),
    .A4(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3436_ (.I(_3172_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3437_ (.A1(\mod.registers.r3[6] ),
    .A2(_3171_),
    .B1(_0464_),
    .B2(\mod.registers.r6[6] ),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3438_ (.A1(\mod.registers.r4[6] ),
    .A2(_3177_),
    .B1(_3181_),
    .B2(\mod.registers.r2[6] ),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3439_ (.I(_3187_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3440_ (.A1(\mod.registers.r7[6] ),
    .A2(_0467_),
    .B1(_3189_),
    .B2(\mod.registers.r12[6] ),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3441_ (.I(_3183_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3442_ (.A1(\mod.registers.r14[6] ),
    .A2(_0469_),
    .B1(_3185_),
    .B2(\mod.registers.r15[6] ),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3443_ (.A1(_0465_),
    .A2(_0466_),
    .A3(_0468_),
    .A4(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3444_ (.A1(_0463_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3445_ (.A1(_0453_),
    .A2(_0456_),
    .B(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3446_ (.I(_3206_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3447_ (.I(_3210_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3448_ (.A1(\mod.registers.r15[6] ),
    .A2(_0474_),
    .B1(_0475_),
    .B2(\mod.registers.r12[6] ),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3449_ (.I(_3225_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3450_ (.I(_3223_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3451_ (.A1(\mod.registers.r2[6] ),
    .A2(_0477_),
    .B1(_0478_),
    .B2(\mod.registers.r3[6] ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3452_ (.I(_3233_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3453_ (.I(_3212_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3454_ (.A1(\mod.registers.r13[6] ),
    .A2(_0480_),
    .B1(_0481_),
    .B2(\mod.registers.r14[6] ),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3455_ (.I(_3230_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3456_ (.I(_3218_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3457_ (.A1(\mod.registers.r1[6] ),
    .A2(_0483_),
    .B1(_0484_),
    .B2(\mod.registers.r4[6] ),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3458_ (.A1(_0476_),
    .A2(_0479_),
    .A3(_0482_),
    .A4(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3459_ (.I(_0422_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3460_ (.I(_0424_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3461_ (.A1(\mod.registers.r5[6] ),
    .A2(_0487_),
    .B1(_0488_),
    .B2(\mod.registers.r9[6] ),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3462_ (.I(_0415_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3463_ (.I(_0417_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3464_ (.A1(\mod.registers.r8[6] ),
    .A2(_0490_),
    .B1(_0491_),
    .B2(\mod.registers.r6[6] ),
    .C1(_0420_),
    .C2(\mod.registers.r11[6] ),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3465_ (.I(_0428_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3466_ (.I(_0430_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3467_ (.A1(\mod.registers.r10[6] ),
    .A2(_0493_),
    .B1(_0494_),
    .B2(\mod.registers.r7[6] ),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3468_ (.A1(_0489_),
    .A2(_0492_),
    .A3(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3469_ (.I(_3195_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3470_ (.A1(_3199_),
    .A2(_0486_),
    .A3(_0496_),
    .B(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3471_ (.I(_3166_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3472_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3473_ (.I(_3232_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3474_ (.I0(\mod.instr_2[4] ),
    .I1(_0501_),
    .S(_0442_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3475_ (.I0(_0502_),
    .I1(\mod.funct3[1] ),
    .S(_0445_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3476_ (.A1(_0500_),
    .A2(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3477_ (.A1(_0473_),
    .A2(_0498_),
    .A3(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3478_ (.I(\mod.pc_2[5] ),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3479_ (.I(_3126_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3480_ (.A1(\mod.registers.r8[5] ),
    .A2(_0457_),
    .B1(_3152_),
    .B2(\mod.registers.r9[5] ),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3481_ (.I(_3143_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3482_ (.A1(\mod.registers.r13[5] ),
    .A2(_3140_),
    .B1(_0509_),
    .B2(\mod.registers.r1[5] ),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3483_ (.A1(\mod.registers.r5[5] ),
    .A2(_0460_),
    .B1(_3160_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3484_ (.A1(\mod.registers.r11[5] ),
    .A2(_3164_),
    .B(_0435_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3485_ (.A1(_0508_),
    .A2(_0510_),
    .A3(_0511_),
    .A4(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3486_ (.A1(\mod.registers.r3[5] ),
    .A2(_3171_),
    .B1(_0464_),
    .B2(\mod.registers.r6[5] ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3487_ (.A1(\mod.registers.r4[5] ),
    .A2(_3177_),
    .B1(_3181_),
    .B2(\mod.registers.r2[5] ),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3488_ (.I(_3189_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3489_ (.A1(\mod.registers.r7[5] ),
    .A2(_0467_),
    .B1(_0516_),
    .B2(\mod.registers.r12[5] ),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3490_ (.I(_3185_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3491_ (.A1(\mod.registers.r14[5] ),
    .A2(_0469_),
    .B1(_0518_),
    .B2(\mod.registers.r15[5] ),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3492_ (.A1(_0514_),
    .A2(_0515_),
    .A3(_0517_),
    .A4(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3493_ (.A1(_0506_),
    .A2(_0507_),
    .B1(_0513_),
    .B2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3494_ (.I(_0499_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3495_ (.I(\mod.instr_2[3] ),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3496_ (.I(_3229_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3497_ (.I0(_0523_),
    .I1(_0524_),
    .S(_0443_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3498_ (.A1(\mod.funct3[0] ),
    .A2(_0439_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3499_ (.A1(_0439_),
    .A2(_0525_),
    .B(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3500_ (.A1(\mod.registers.r13[5] ),
    .A2(_3234_),
    .B1(_3213_),
    .B2(\mod.registers.r14[5] ),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3501_ (.A1(\mod.registers.r8[5] ),
    .A2(_0416_),
    .B1(_0420_),
    .B2(\mod.registers.r11[5] ),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3502_ (.A1(\mod.registers.r15[5] ),
    .A2(_0474_),
    .B1(_0475_),
    .B2(\mod.registers.r12[5] ),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3503_ (.A1(\mod.registers.r9[5] ),
    .A2(_0425_),
    .B1(_0429_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3504_ (.A1(_0528_),
    .A2(_0529_),
    .A3(_0530_),
    .A4(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3505_ (.A1(\mod.registers.r7[5] ),
    .A2(_0431_),
    .B1(_3224_),
    .B2(\mod.registers.r3[5] ),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3506_ (.A1(\mod.registers.r5[5] ),
    .A2(_0423_),
    .B1(_3219_),
    .B2(\mod.registers.r4[5] ),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3507_ (.A1(\mod.registers.r6[5] ),
    .A2(_0417_),
    .B1(_3226_),
    .B2(\mod.registers.r2[5] ),
    .C1(_3230_),
    .C2(\mod.registers.r1[5] ),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3508_ (.A1(_0533_),
    .A2(_0534_),
    .A3(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3509_ (.A1(_0532_),
    .A2(_0536_),
    .B(_3108_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(_3107_),
    .A2(_3165_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3511_ (.I(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3512_ (.I(\mod.funct7[1] ),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3513_ (.I0(_3194_),
    .I1(_0540_),
    .S(_0443_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3514_ (.A1(_0539_),
    .A2(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3515_ (.A1(_0522_),
    .A2(_0527_),
    .B(_0537_),
    .C(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3516_ (.A1(_0521_),
    .A2(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3517_ (.I(_0500_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3518_ (.I(_3198_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3519_ (.I(_0428_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3520_ (.I(_0419_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3521_ (.A1(\mod.registers.r10[4] ),
    .A2(_0547_),
    .B1(_0548_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3522_ (.A1(\mod.registers.r2[4] ),
    .A2(_0477_),
    .B1(_0488_),
    .B2(\mod.registers.r9[4] ),
    .C1(\mod.registers.r13[4] ),
    .C2(_0480_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3523_ (.I(_0430_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3524_ (.A1(\mod.registers.r1[4] ),
    .A2(_0483_),
    .B1(_0551_),
    .B2(\mod.registers.r7[4] ),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3525_ (.A1(_0549_),
    .A2(_0550_),
    .A3(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3526_ (.A1(\mod.registers.r14[4] ),
    .A2(_0481_),
    .B1(_0478_),
    .B2(\mod.registers.r3[4] ),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3527_ (.I(_3210_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3528_ (.A1(\mod.registers.r8[4] ),
    .A2(_0490_),
    .B1(_0555_),
    .B2(\mod.registers.r12[4] ),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3529_ (.A1(\mod.registers.r6[4] ),
    .A2(_0491_),
    .B1(_0484_),
    .B2(\mod.registers.r4[4] ),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3530_ (.I(_3206_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3531_ (.I(_0422_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3532_ (.A1(\mod.registers.r15[4] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\mod.registers.r5[4] ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3533_ (.A1(_0554_),
    .A2(_0556_),
    .A3(_0557_),
    .A4(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3534_ (.I(_3198_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3535_ (.I(\mod.funct7[0] ),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3536_ (.I0(_0540_),
    .I1(_0563_),
    .S(_0443_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3537_ (.A1(_0562_),
    .A2(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3538_ (.A1(_0546_),
    .A2(_0553_),
    .A3(_0561_),
    .B(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3539_ (.A1(_0545_),
    .A2(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3540_ (.I(\mod.pc_2[4] ),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3541_ (.I(_0436_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3542_ (.I(_3176_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3543_ (.I(_3180_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3544_ (.I(_3172_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3545_ (.A1(\mod.registers.r4[4] ),
    .A2(_0570_),
    .B1(_0571_),
    .B2(\mod.registers.r2[4] ),
    .C1(_0572_),
    .C2(\mod.registers.r6[4] ),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3546_ (.A1(\mod.registers.r15[4] ),
    .A2(_0518_),
    .B1(_0509_),
    .B2(\mod.registers.r1[4] ),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3547_ (.A1(\mod.registers.r14[4] ),
    .A2(_0469_),
    .B1(_3164_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3548_ (.I(_3139_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3549_ (.A1(\mod.registers.r9[4] ),
    .A2(_3152_),
    .B1(_0576_),
    .B2(\mod.registers.r13[4] ),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3550_ (.I(_3159_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3551_ (.A1(\mod.registers.r10[4] ),
    .A2(_0578_),
    .B(_0435_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3552_ (.A1(_0574_),
    .A2(_0575_),
    .A3(_0577_),
    .A4(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3553_ (.I(_3150_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3554_ (.I(_3170_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3555_ (.I(_3156_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3556_ (.A1(\mod.registers.r8[4] ),
    .A2(_0581_),
    .B1(_0582_),
    .B2(\mod.registers.r3[4] ),
    .C1(_0583_),
    .C2(\mod.registers.r5[4] ),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3557_ (.I(_0467_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3558_ (.I(_3189_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3559_ (.A1(\mod.registers.r7[4] ),
    .A2(_0585_),
    .B1(_0586_),
    .B2(\mod.registers.r12[4] ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3560_ (.A1(_0573_),
    .A2(_0580_),
    .A3(_0584_),
    .A4(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3561_ (.A1(_0568_),
    .A2(_0569_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3562_ (.A1(_0567_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3563_ (.I(\mod.pc_2[5] ),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3564_ (.A1(_0513_),
    .A2(_0520_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3565_ (.A1(_0591_),
    .A2(_0455_),
    .B(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3566_ (.A1(_0593_),
    .A2(_0543_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3567_ (.A1(_0544_),
    .A2(_0590_),
    .B(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3568_ (.I(\mod.pc_2[7] ),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3569_ (.A1(_0596_),
    .A2(_0436_),
    .B1(_3169_),
    .B2(_3191_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3570_ (.A1(_0597_),
    .A2(_0449_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3571_ (.A1(\mod.pc_2[6] ),
    .A2(_3126_),
    .B1(_0463_),
    .B2(_0471_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3572_ (.A1(_0498_),
    .A2(_0504_),
    .B(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3573_ (.A1(_0599_),
    .A2(_0498_),
    .A3(_0504_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3574_ (.A1(_0600_),
    .A2(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3575_ (.A1(_0598_),
    .A2(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3576_ (.A1(_3193_),
    .A2(_0450_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3577_ (.A1(_0451_),
    .A2(_0505_),
    .B1(_0595_),
    .B2(_0603_),
    .C(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3578_ (.A1(\mod.registers.r7[2] ),
    .A2(_0494_),
    .B1(_0478_),
    .B2(\mod.registers.r3[2] ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3579_ (.A1(\mod.registers.r1[2] ),
    .A2(_0483_),
    .B1(_0484_),
    .B2(\mod.registers.r4[2] ),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3580_ (.A1(_0606_),
    .A2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3581_ (.A1(\mod.registers.r5[2] ),
    .A2(_0423_),
    .B1(_3226_),
    .B2(\mod.registers.r2[2] ),
    .C1(_0491_),
    .C2(\mod.registers.r6[2] ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3582_ (.A1(\mod.registers.r9[2] ),
    .A2(_0488_),
    .B1(_0493_),
    .B2(\mod.registers.r10[2] ),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3583_ (.A1(\mod.registers.r8[2] ),
    .A2(_0490_),
    .B1(_0548_),
    .B2(\mod.registers.r11[2] ),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3584_ (.I(\mod.registers.r12[2] ),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3585_ (.I(_3209_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3586_ (.A1(_3215_),
    .A2(_0414_),
    .A3(_3232_),
    .A4(_3205_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3587_ (.I(\mod.registers.r15[2] ),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3588_ (.A1(_0612_),
    .A2(_3208_),
    .A3(_0613_),
    .B1(_0614_),
    .B2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3589_ (.A1(\mod.registers.r13[2] ),
    .A2(_0480_),
    .B1(_0481_),
    .B2(\mod.registers.r14[2] ),
    .C(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3590_ (.A1(_0609_),
    .A2(_0610_),
    .A3(_0611_),
    .A4(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3591_ (.A1(_0546_),
    .A2(_0608_),
    .A3(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3592_ (.A1(_3108_),
    .A2(_0444_),
    .B(_0500_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3593_ (.A1(_0619_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3594_ (.I(\mod.pc_2[2] ),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3595_ (.A1(\mod.registers.r8[2] ),
    .A2(_0457_),
    .B1(_3160_),
    .B2(\mod.registers.r10[2] ),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3596_ (.I(_3183_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3597_ (.A1(\mod.registers.r14[2] ),
    .A2(_0624_),
    .B1(_0464_),
    .B2(\mod.registers.r6[2] ),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3598_ (.I(_3163_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3599_ (.A1(\mod.registers.r11[2] ),
    .A2(_0626_),
    .B1(_0571_),
    .B2(\mod.registers.r2[2] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3600_ (.I(_3176_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3601_ (.A1(\mod.registers.r4[2] ),
    .A2(_0628_),
    .B(_0499_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3602_ (.A1(_0623_),
    .A2(_0625_),
    .A3(_0627_),
    .A4(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3603_ (.A1(\mod.registers.r5[2] ),
    .A2(_0583_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3604_ (.I(_3187_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3605_ (.A1(\mod.registers.r7[2] ),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3606_ (.I(_3175_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3607_ (.I(_3137_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3608_ (.A1(_3174_),
    .A2(_0635_),
    .A3(_3134_),
    .A4(_3179_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3609_ (.A1(_0612_),
    .A2(_0634_),
    .A3(_3188_),
    .B1(_0636_),
    .B2(_0615_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3610_ (.A1(\mod.registers.r13[2] ),
    .A2(_3140_),
    .B1(_3144_),
    .B2(\mod.registers.r1[2] ),
    .C(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3611_ (.I(_3151_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3612_ (.A1(\mod.registers.r9[2] ),
    .A2(_0639_),
    .B1(_0582_),
    .B2(\mod.registers.r3[2] ),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3613_ (.A1(_0631_),
    .A2(_0633_),
    .A3(_0638_),
    .A4(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3614_ (.A1(_0622_),
    .A2(_0522_),
    .B1(_0630_),
    .B2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3615_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3616_ (.A1(_0621_),
    .A2(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3617_ (.I(_3198_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3618_ (.A1(\mod.registers.r7[3] ),
    .A2(_0431_),
    .B1(_3224_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3619_ (.A1(\mod.registers.r1[3] ),
    .A2(_3231_),
    .B1(_3219_),
    .B2(\mod.registers.r4[3] ),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_0646_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3621_ (.A1(\mod.registers.r5[3] ),
    .A2(_0423_),
    .B1(_3226_),
    .B2(\mod.registers.r2[3] ),
    .C1(_0418_),
    .C2(\mod.registers.r6[3] ),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3622_ (.A1(\mod.registers.r9[3] ),
    .A2(_0425_),
    .B1(_0429_),
    .B2(\mod.registers.r10[3] ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3623_ (.A1(\mod.registers.r8[3] ),
    .A2(_0416_),
    .B1(_0420_),
    .B2(\mod.registers.r11[3] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3624_ (.I(\mod.registers.r12[3] ),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3625_ (.I(\mod.registers.r15[3] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3626_ (.A1(_0652_),
    .A2(_3208_),
    .A3(_0613_),
    .B1(_0614_),
    .B2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3627_ (.A1(\mod.registers.r13[3] ),
    .A2(_3234_),
    .B1(_3213_),
    .B2(\mod.registers.r14[3] ),
    .C(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3628_ (.A1(_0649_),
    .A2(_0650_),
    .A3(_0651_),
    .A4(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3629_ (.I(_3215_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3630_ (.I0(\mod.funct7[0] ),
    .I1(_0657_),
    .S(_0442_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3631_ (.A1(_0538_),
    .A2(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3632_ (.A1(_0645_),
    .A2(_0648_),
    .A3(_0656_),
    .B(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3633_ (.I(_3126_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3634_ (.A1(\mod.registers.r8[3] ),
    .A2(_3150_),
    .B1(_3159_),
    .B2(\mod.registers.r10[3] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3635_ (.A1(\mod.registers.r14[3] ),
    .A2(_3183_),
    .B1(_3172_),
    .B2(\mod.registers.r6[3] ),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3636_ (.A1(\mod.registers.r11[3] ),
    .A2(_3163_),
    .B1(_3180_),
    .B2(\mod.registers.r2[3] ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3637_ (.A1(\mod.registers.r4[3] ),
    .A2(_3177_),
    .B(_3167_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3638_ (.A1(_0662_),
    .A2(_0663_),
    .A3(_0664_),
    .A4(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3639_ (.A1(\mod.registers.r5[3] ),
    .A2(_0460_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3640_ (.A1(\mod.registers.r7[3] ),
    .A2(_3187_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3641_ (.A1(\mod.registers.r9[3] ),
    .A2(_3151_),
    .B1(_3170_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3642_ (.A1(_0652_),
    .A2(_3175_),
    .A3(_3188_),
    .B1(_0636_),
    .B2(_0653_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3643_ (.A1(\mod.registers.r13[3] ),
    .A2(_3139_),
    .B1(_3143_),
    .B2(\mod.registers.r1[3] ),
    .C(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3644_ (.A1(_0667_),
    .A2(_0668_),
    .A3(_0669_),
    .A4(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3645_ (.A1(\mod.pc_2[3] ),
    .A2(_0661_),
    .B1(_0666_),
    .B2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3646_ (.A1(_0455_),
    .A2(_0660_),
    .A3(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3647_ (.A1(_0648_),
    .A2(_0656_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3648_ (.I(\mod.pc_2[3] ),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(_0435_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3650_ (.A1(_0662_),
    .A2(_0663_),
    .A3(_0664_),
    .A4(_0665_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3651_ (.A1(_0667_),
    .A2(_0668_),
    .A3(_0669_),
    .A4(_0671_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3652_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0678_),
    .B2(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3653_ (.A1(_0546_),
    .A2(_0658_),
    .B1(_0675_),
    .B2(_3106_),
    .C(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3654_ (.A1(_0674_),
    .A2(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3655_ (.A1(_0456_),
    .A2(_0660_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3656_ (.I(_0680_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3657_ (.A1(_0683_),
    .A2(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3658_ (.A1(_0644_),
    .A2(_0682_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3659_ (.A1(\mod.registers.r1[1] ),
    .A2(_3231_),
    .B1(_3219_),
    .B2(\mod.registers.r4[1] ),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3660_ (.A1(\mod.registers.r5[1] ),
    .A2(_0487_),
    .B1(_0477_),
    .B2(\mod.registers.r2[1] ),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3661_ (.A1(_0687_),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3662_ (.A1(\mod.registers.r6[1] ),
    .A2(_0418_),
    .B1(_3223_),
    .B2(\mod.registers.r3[1] ),
    .C1(_0430_),
    .C2(\mod.registers.r7[1] ),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3663_ (.A1(\mod.registers.r8[1] ),
    .A2(_0416_),
    .B1(_0425_),
    .B2(\mod.registers.r9[1] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3664_ (.A1(\mod.registers.r10[1] ),
    .A2(_0429_),
    .B1(_0548_),
    .B2(\mod.registers.r11[1] ),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3665_ (.I(_3202_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3666_ (.A1(_3215_),
    .A2(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3667_ (.I(_3220_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3668_ (.A1(_3232_),
    .A2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3669_ (.A1(\mod.registers.r12[1] ),
    .A2(_0694_),
    .A3(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3670_ (.A1(_0501_),
    .A2(_0524_),
    .A3(\mod.registers.r14[1] ),
    .A4(_0694_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3671_ (.A1(_0427_),
    .A2(_0695_),
    .A3(\mod.registers.r13[1] ),
    .A4(_0694_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3672_ (.A1(\mod.registers.r15[1] ),
    .A2(_3206_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3673_ (.A1(_0697_),
    .A2(_0698_),
    .A3(_0699_),
    .A4(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3674_ (.A1(_0690_),
    .A2(_0691_),
    .A3(_0692_),
    .A4(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3675_ (.A1(_0562_),
    .A2(_0689_),
    .A3(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3676_ (.A1(_3106_),
    .A2(_0502_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3677_ (.A1(_0522_),
    .A2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3678_ (.A1(_0703_),
    .A2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3679_ (.I(\mod.pc_2[1] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3680_ (.A1(\mod.registers.r8[1] ),
    .A2(_0581_),
    .B1(_0576_),
    .B2(\mod.registers.r13[1] ),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3681_ (.A1(\mod.registers.r6[1] ),
    .A2(_0572_),
    .B1(_0516_),
    .B2(\mod.registers.r12[1] ),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(_3179_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3683_ (.I(_3174_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3684_ (.A1(_0711_),
    .A2(_0635_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3685_ (.A1(_3178_),
    .A2(_0710_),
    .A3(\mod.registers.r1[1] ),
    .A4(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3686_ (.I(_3134_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3687_ (.A1(_0714_),
    .A2(_0710_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3688_ (.A1(_3147_),
    .A2(_0635_),
    .A3(\mod.registers.r4[1] ),
    .A4(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3689_ (.A1(_0714_),
    .A2(_3136_),
    .A3(\mod.registers.r2[1] ),
    .A4(_0712_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3690_ (.A1(_3125_),
    .A2(_0713_),
    .A3(_0716_),
    .A4(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3691_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3692_ (.A1(\mod.registers.r15[1] ),
    .A2(_0518_),
    .B1(_0582_),
    .B2(\mod.registers.r3[1] ),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3693_ (.A1(\mod.registers.r14[1] ),
    .A2(_0624_),
    .B1(_0626_),
    .B2(\mod.registers.r11[1] ),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3694_ (.A1(\mod.registers.r9[1] ),
    .A2(_0639_),
    .B1(_0578_),
    .B2(\mod.registers.r10[1] ),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3695_ (.A1(\mod.registers.r7[1] ),
    .A2(_0632_),
    .B1(_0583_),
    .B2(\mod.registers.r5[1] ),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3696_ (.A1(_0720_),
    .A2(_0721_),
    .A3(_0722_),
    .A4(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3697_ (.A1(_0707_),
    .A2(_0455_),
    .B1(_0719_),
    .B2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3698_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3699_ (.A1(_0706_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3700_ (.A1(_0539_),
    .A2(_0502_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3701_ (.A1(_3199_),
    .A2(_0689_),
    .A3(_0702_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3702_ (.I(\mod.pc_2[1] ),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3703_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0718_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3704_ (.A1(_0720_),
    .A2(_0721_),
    .A3(_0722_),
    .A4(_0723_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3705_ (.A1(_0730_),
    .A2(_0507_),
    .B1(_0731_),
    .B2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3706_ (.A1(_0545_),
    .A2(_0729_),
    .A3(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3707_ (.A1(_0703_),
    .A2(_0705_),
    .B(_0725_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3708_ (.A1(\mod.registers.r7[0] ),
    .A2(_0431_),
    .B1(_3224_),
    .B2(\mod.registers.r3[0] ),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3709_ (.A1(\mod.registers.r1[0] ),
    .A2(_3231_),
    .B1(_3218_),
    .B2(\mod.registers.r4[0] ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3710_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3711_ (.A1(\mod.registers.r5[0] ),
    .A2(_0422_),
    .B1(_3225_),
    .B2(\mod.registers.r2[0] ),
    .C1(_0417_),
    .C2(\mod.registers.r6[0] ),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3712_ (.A1(\mod.registers.r9[0] ),
    .A2(_0424_),
    .B1(_0428_),
    .B2(\mod.registers.r10[0] ),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3713_ (.A1(\mod.registers.r8[0] ),
    .A2(_0415_),
    .B1(_0419_),
    .B2(\mod.registers.r11[0] ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3714_ (.I(\mod.registers.r12[0] ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3715_ (.I(\mod.registers.r15[0] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3716_ (.A1(_0742_),
    .A2(_3208_),
    .A3(_0613_),
    .B1(_0614_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3717_ (.A1(\mod.registers.r13[0] ),
    .A2(_3233_),
    .B1(_3212_),
    .B2(\mod.registers.r14[0] ),
    .C(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3718_ (.A1(_0739_),
    .A2(_0740_),
    .A3(_0741_),
    .A4(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3719_ (.A1(_0645_),
    .A2(_0738_),
    .A3(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3720_ (.A1(_3108_),
    .A2(_0525_),
    .B(_0454_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3721_ (.A1(\mod.registers.r8[0] ),
    .A2(_0581_),
    .B1(_0578_),
    .B2(\mod.registers.r10[0] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3722_ (.A1(\mod.registers.r14[0] ),
    .A2(_0624_),
    .B1(_0572_),
    .B2(\mod.registers.r6[0] ),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3723_ (.A1(\mod.registers.r11[0] ),
    .A2(_0626_),
    .B1(_0571_),
    .B2(\mod.registers.r2[0] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3724_ (.A1(\mod.registers.r4[0] ),
    .A2(_0628_),
    .B(_0499_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3725_ (.A1(_0749_),
    .A2(_0750_),
    .A3(_0751_),
    .A4(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3726_ (.A1(\mod.registers.r7[0] ),
    .A2(_0632_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3727_ (.A1(\mod.registers.r5[0] ),
    .A2(_0583_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3728_ (.A1(_0742_),
    .A2(_0634_),
    .A3(_3188_),
    .B1(_0636_),
    .B2(_0743_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3729_ (.A1(\mod.registers.r13[0] ),
    .A2(_0576_),
    .B1(_0509_),
    .B2(\mod.registers.r1[0] ),
    .C(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3730_ (.A1(\mod.registers.r9[0] ),
    .A2(_0639_),
    .B1(_0582_),
    .B2(\mod.registers.r3[0] ),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3731_ (.A1(_0754_),
    .A2(_0755_),
    .A3(_0757_),
    .A4(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3732_ (.A1(\mod.pc_2[0] ),
    .A2(_0507_),
    .B1(_0753_),
    .B2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3733_ (.A1(_0747_),
    .A2(_0748_),
    .A3(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3734_ (.A1(_0734_),
    .A2(_0735_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3735_ (.I(_0677_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3736_ (.A1(_3199_),
    .A2(_0444_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3737_ (.A1(_0562_),
    .A2(_0608_),
    .A3(_0618_),
    .B(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3738_ (.I(\mod.pc_2[2] ),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3739_ (.A1(_0623_),
    .A2(_0625_),
    .A3(_0627_),
    .A4(_0629_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3740_ (.A1(_0631_),
    .A2(_0633_),
    .A3(_0638_),
    .A4(_0640_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3741_ (.A1(_0766_),
    .A2(_0661_),
    .B1(_0767_),
    .B2(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3742_ (.A1(_0763_),
    .A2(_0765_),
    .A3(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3743_ (.A1(_0619_),
    .A2(_0620_),
    .B(_0642_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3744_ (.A1(_0770_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3745_ (.A1(_0727_),
    .A2(_0762_),
    .B(_0772_),
    .C(_0682_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3746_ (.A1(_0598_),
    .A2(_0602_),
    .A3(_0544_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3747_ (.A1(_0545_),
    .A2(_0566_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3748_ (.A1(_0763_),
    .A2(_0566_),
    .A3(_0588_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3749_ (.A1(_0775_),
    .A2(_0589_),
    .B(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3750_ (.A1(_0686_),
    .A2(_0773_),
    .B(_0774_),
    .C(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3751_ (.I(\mod.pc_2[8] ),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3752_ (.I(_0500_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3753_ (.I(_3151_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3754_ (.I(_3170_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3755_ (.A1(\mod.registers.r9[8] ),
    .A2(_0781_),
    .B1(_0782_),
    .B2(\mod.registers.r3[8] ),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3756_ (.I(_3139_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3757_ (.A1(\mod.registers.r13[8] ),
    .A2(_0784_),
    .B1(_0586_),
    .B2(\mod.registers.r12[8] ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3758_ (.I(_3156_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3759_ (.A1(\mod.registers.r5[8] ),
    .A2(_0786_),
    .B(_0677_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3760_ (.I(_3185_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3761_ (.A1(\mod.registers.r7[8] ),
    .A2(_0585_),
    .B1(_0788_),
    .B2(\mod.registers.r15[8] ),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3762_ (.A1(_0783_),
    .A2(_0785_),
    .A3(_0787_),
    .A4(_0789_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3763_ (.I(_0457_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3764_ (.I(_3181_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3765_ (.A1(\mod.registers.r8[8] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\mod.registers.r2[8] ),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_3144_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3767_ (.A1(\mod.registers.r4[8] ),
    .A2(_0570_),
    .B1(_0794_),
    .B2(\mod.registers.r1[8] ),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3768_ (.I(_0469_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3769_ (.I(_3159_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3770_ (.A1(\mod.registers.r14[8] ),
    .A2(_0796_),
    .B1(_0797_),
    .B2(\mod.registers.r10[8] ),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3771_ (.I(_3163_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3772_ (.I(_0464_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3773_ (.A1(\mod.registers.r11[8] ),
    .A2(_0799_),
    .B1(_0800_),
    .B2(\mod.registers.r6[8] ),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3774_ (.A1(_0793_),
    .A2(_0795_),
    .A3(_0798_),
    .A4(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3775_ (.A1(_0779_),
    .A2(_0780_),
    .B1(_0790_),
    .B2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3776_ (.I(_0645_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3777_ (.I(_0488_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3778_ (.I(_3218_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3779_ (.A1(\mod.registers.r9[8] ),
    .A2(_0805_),
    .B1(_0806_),
    .B2(\mod.registers.r4[8] ),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3780_ (.I(_0419_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3781_ (.A1(\mod.registers.r10[8] ),
    .A2(_0547_),
    .B1(_0808_),
    .B2(\mod.registers.r11[8] ),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3782_ (.I(_0474_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3783_ (.I(_0478_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3784_ (.A1(\mod.registers.r15[8] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(\mod.registers.r3[8] ),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3785_ (.I(_0490_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3786_ (.A1(\mod.registers.r8[8] ),
    .A2(_0813_),
    .B1(_0551_),
    .B2(\mod.registers.r7[8] ),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3787_ (.A1(_0807_),
    .A2(_0809_),
    .A3(_0812_),
    .A4(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3788_ (.I(_0418_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3789_ (.I(_3234_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3790_ (.A1(\mod.registers.r6[8] ),
    .A2(_0816_),
    .B1(_0555_),
    .B2(\mod.registers.r12[8] ),
    .C1(\mod.registers.r13[8] ),
    .C2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3791_ (.I(_0487_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3792_ (.I(_3213_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3793_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3794_ (.A1(\mod.registers.r5[8] ),
    .A2(_0819_),
    .B1(_0821_),
    .B2(\mod.registers.r14[8] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3795_ (.I(_0477_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3796_ (.I(_0483_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3797_ (.A1(\mod.registers.r2[8] ),
    .A2(_0823_),
    .B1(_0824_),
    .B2(\mod.registers.r1[8] ),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3798_ (.A1(_0818_),
    .A2(_0822_),
    .A3(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3799_ (.I(_0497_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3800_ (.A1(_0804_),
    .A2(_0815_),
    .A3(_0826_),
    .B(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3801_ (.I(_0445_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3802_ (.I0(_0658_),
    .I1(_0710_),
    .S(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3803_ (.A1(_0456_),
    .A2(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3804_ (.A1(_0803_),
    .A2(_0828_),
    .A3(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3805_ (.I(\mod.pc_2[8] ),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3806_ (.I(_0507_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3807_ (.A1(_0783_),
    .A2(_0785_),
    .A3(_0787_),
    .A4(_0789_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3808_ (.A1(_0793_),
    .A2(_0795_),
    .A3(_0798_),
    .A4(_0801_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3809_ (.A1(_0833_),
    .A2(_0834_),
    .B1(_0835_),
    .B2(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(_0828_),
    .A2(_0831_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3811_ (.A1(_0837_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(_0832_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3813_ (.A1(\mod.pc_2[9] ),
    .A2(_0661_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3814_ (.A1(\mod.registers.r14[9] ),
    .A2(_0796_),
    .B1(_0800_),
    .B2(\mod.registers.r6[9] ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3815_ (.A1(\mod.registers.r1[9] ),
    .A2(_0794_),
    .B1(_0792_),
    .B2(\mod.registers.r2[9] ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3816_ (.A1(_0842_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3817_ (.A1(\mod.registers.r8[9] ),
    .A2(_0791_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3818_ (.A1(\mod.registers.r3[9] ),
    .A2(_0782_),
    .B1(_0797_),
    .B2(\mod.registers.r10[9] ),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3819_ (.A1(_0661_),
    .A2(_0845_),
    .A3(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3820_ (.A1(\mod.registers.r11[9] ),
    .A2(_0799_),
    .B1(_0786_),
    .B2(\mod.registers.r5[9] ),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3821_ (.A1(\mod.registers.r7[9] ),
    .A2(_0632_),
    .B1(_0788_),
    .B2(\mod.registers.r15[9] ),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3822_ (.A1(\mod.registers.r4[9] ),
    .A2(_0628_),
    .B1(_0784_),
    .B2(\mod.registers.r13[9] ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3823_ (.A1(\mod.registers.r9[9] ),
    .A2(_0781_),
    .B1(_0516_),
    .B2(\mod.registers.r12[9] ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3824_ (.A1(_0848_),
    .A2(_0849_),
    .A3(_0850_),
    .A4(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3825_ (.A1(_0844_),
    .A2(_0847_),
    .A3(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3826_ (.A1(_0841_),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3827_ (.I(_0424_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3828_ (.A1(\mod.registers.r5[9] ),
    .A2(_0559_),
    .B1(_0806_),
    .B2(\mod.registers.r4[9] ),
    .C1(_0855_),
    .C2(\mod.registers.r9[9] ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3829_ (.A1(\mod.registers.r15[9] ),
    .A2(_0558_),
    .B1(_0555_),
    .B2(\mod.registers.r12[9] ),
    .C1(_0551_),
    .C2(\mod.registers.r7[9] ),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3830_ (.I(_0415_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_3223_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3832_ (.A1(\mod.registers.r8[9] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\mod.registers.r3[9] ),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3833_ (.A1(_0856_),
    .A2(_0857_),
    .A3(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3834_ (.A1(\mod.registers.r13[9] ),
    .A2(_0817_),
    .B1(_0808_),
    .B2(\mod.registers.r11[9] ),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3835_ (.I(_3230_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3836_ (.A1(\mod.registers.r6[9] ),
    .A2(_0816_),
    .B1(_0863_),
    .B2(\mod.registers.r1[9] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3837_ (.I(_3225_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3838_ (.A1(\mod.registers.r2[9] ),
    .A2(_0865_),
    .B1(_0547_),
    .B2(\mod.registers.r10[9] ),
    .C1(\mod.registers.r14[9] ),
    .C2(_0820_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3839_ (.A1(_0862_),
    .A2(_0864_),
    .A3(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3840_ (.A1(_0804_),
    .A2(_0861_),
    .A3(_0867_),
    .B(_0497_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_0445_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(_0714_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3843_ (.A1(_0869_),
    .A2(_0564_),
    .B(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3844_ (.A1(_0763_),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3845_ (.A1(_0868_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(_0854_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3847_ (.A1(_0841_),
    .A2(_0853_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3848_ (.A1(_0875_),
    .A2(_0868_),
    .A3(_0872_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3849_ (.A1(_0874_),
    .A2(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3850_ (.I(\mod.pc_2[11] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3851_ (.A1(\mod.registers.r8[11] ),
    .A2(_0791_),
    .B1(_0797_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3852_ (.A1(\mod.registers.r13[11] ),
    .A2(_0784_),
    .B1(_0788_),
    .B2(\mod.registers.r15[11] ),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3853_ (.A1(\mod.registers.r14[11] ),
    .A2(_0796_),
    .B(_0454_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3854_ (.A1(\mod.registers.r3[11] ),
    .A2(_0782_),
    .B1(_0800_),
    .B2(\mod.registers.r6[11] ),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3855_ (.A1(_0879_),
    .A2(_0880_),
    .A3(_0881_),
    .A4(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3856_ (.A1(\mod.registers.r9[11] ),
    .A2(_0781_),
    .B1(_0794_),
    .B2(\mod.registers.r1[11] ),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3857_ (.A1(\mod.registers.r7[11] ),
    .A2(_0585_),
    .B1(_0586_),
    .B2(\mod.registers.r12[11] ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3858_ (.A1(\mod.registers.r4[11] ),
    .A2(_0570_),
    .B1(_0799_),
    .B2(\mod.registers.r11[11] ),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3859_ (.A1(\mod.registers.r5[11] ),
    .A2(_0786_),
    .B1(_0792_),
    .B2(\mod.registers.r2[11] ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3860_ (.A1(_0884_),
    .A2(_0885_),
    .A3(_0886_),
    .A4(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3861_ (.A1(_0883_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3862_ (.A1(_0878_),
    .A2(_0780_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3863_ (.A1(\mod.registers.r15[11] ),
    .A2(_0558_),
    .B1(_0551_),
    .B2(\mod.registers.r7[11] ),
    .C1(_0859_),
    .C2(\mod.registers.r3[11] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3864_ (.A1(\mod.registers.r5[11] ),
    .A2(_0559_),
    .B1(_0806_),
    .B2(\mod.registers.r4[11] ),
    .C1(_0858_),
    .C2(\mod.registers.r8[11] ),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3865_ (.I(_0475_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3866_ (.A1(\mod.registers.r12[11] ),
    .A2(_0893_),
    .B1(_0547_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3867_ (.A1(_0891_),
    .A2(_0892_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3868_ (.A1(\mod.registers.r2[11] ),
    .A2(_0865_),
    .B1(_0855_),
    .B2(\mod.registers.r9[11] ),
    .C1(\mod.registers.r14[11] ),
    .C2(_0820_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3869_ (.A1(\mod.registers.r1[11] ),
    .A2(_0863_),
    .B1(_0808_),
    .B2(\mod.registers.r11[11] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3870_ (.I(_0491_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3871_ (.A1(\mod.registers.r6[11] ),
    .A2(_0898_),
    .B1(_0817_),
    .B2(\mod.registers.r13[11] ),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3872_ (.A1(_0896_),
    .A2(_0897_),
    .A3(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3873_ (.A1(_0804_),
    .A2(_0895_),
    .A3(_0900_),
    .B(_0827_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3874_ (.A1(\mod.funct7[2] ),
    .A2(_0869_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3875_ (.A1(_3147_),
    .A2(_0829_),
    .B(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3876_ (.A1(_0545_),
    .A2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3877_ (.A1(_0901_),
    .A2(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3878_ (.A1(_0890_),
    .A2(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_0878_),
    .A2(_0763_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3880_ (.A1(_0883_),
    .A2(_0888_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3881_ (.A1(_0908_),
    .A2(_0901_),
    .A3(_0904_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_0906_),
    .A2(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3883_ (.I(\mod.pc_2[10] ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3884_ (.A1(\mod.registers.r14[10] ),
    .A2(_0796_),
    .B1(_0786_),
    .B2(\mod.registers.r5[10] ),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3885_ (.A1(\mod.registers.r6[10] ),
    .A2(_0800_),
    .B1(_0792_),
    .B2(\mod.registers.r2[10] ),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3886_ (.A1(\mod.registers.r13[10] ),
    .A2(_0784_),
    .B1(_0794_),
    .B2(\mod.registers.r1[10] ),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3887_ (.A1(\mod.registers.r7[10] ),
    .A2(_0585_),
    .B(_0677_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3888_ (.A1(_0912_),
    .A2(_0913_),
    .A3(_0914_),
    .A4(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3889_ (.A1(\mod.registers.r9[10] ),
    .A2(_0781_),
    .B1(_0788_),
    .B2(\mod.registers.r15[10] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3890_ (.A1(\mod.registers.r3[10] ),
    .A2(_0782_),
    .B1(_0586_),
    .B2(\mod.registers.r12[10] ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3891_ (.A1(\mod.registers.r8[10] ),
    .A2(_0791_),
    .B1(_0797_),
    .B2(\mod.registers.r10[10] ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3892_ (.A1(\mod.registers.r4[10] ),
    .A2(_0570_),
    .B1(_0799_),
    .B2(\mod.registers.r11[10] ),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3893_ (.A1(_0917_),
    .A2(_0918_),
    .A3(_0919_),
    .A4(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3894_ (.A1(_0911_),
    .A2(_0569_),
    .B1(_0916_),
    .B2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3895_ (.A1(\mod.registers.r8[10] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\mod.registers.r3[10] ),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3896_ (.A1(\mod.registers.r15[10] ),
    .A2(_0474_),
    .B1(_0493_),
    .B2(\mod.registers.r10[10] ),
    .C1(_0494_),
    .C2(\mod.registers.r7[10] ),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3897_ (.A1(\mod.registers.r5[10] ),
    .A2(_0487_),
    .B1(_0484_),
    .B2(\mod.registers.r4[10] ),
    .C1(_0475_),
    .C2(\mod.registers.r12[10] ),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3898_ (.A1(_0923_),
    .A2(_0924_),
    .A3(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3899_ (.A1(\mod.registers.r6[10] ),
    .A2(_0816_),
    .B1(_0817_),
    .B2(\mod.registers.r13[10] ),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3900_ (.A1(\mod.registers.r1[10] ),
    .A2(_0863_),
    .B1(_0808_),
    .B2(\mod.registers.r11[10] ),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3901_ (.A1(\mod.registers.r2[10] ),
    .A2(_0865_),
    .B1(_0855_),
    .B2(\mod.registers.r9[10] ),
    .C1(\mod.registers.r14[10] ),
    .C2(_0481_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3902_ (.A1(_0927_),
    .A2(_0928_),
    .A3(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3903_ (.A1(_0546_),
    .A2(_0926_),
    .A3(_0930_),
    .B(_0497_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3904_ (.I(_0454_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3905_ (.I(_0635_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3906_ (.A1(_0933_),
    .A2(_0439_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3907_ (.A1(_0869_),
    .A2(_0541_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3908_ (.A1(_0932_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3909_ (.A1(_0931_),
    .A2(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3910_ (.A1(_0922_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3911_ (.A1(_0912_),
    .A2(_0913_),
    .A3(_0914_),
    .A4(_0915_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3912_ (.A1(_0917_),
    .A2(_0918_),
    .A3(_0919_),
    .A4(_0920_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3913_ (.A1(\mod.pc_2[10] ),
    .A2(_3127_),
    .B1(_0939_),
    .B2(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3914_ (.A1(_0941_),
    .A2(_0931_),
    .A3(_0936_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3915_ (.A1(_0938_),
    .A2(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3916_ (.A1(_0877_),
    .A2(_0910_),
    .A3(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3917_ (.A1(_0605_),
    .A2(_0778_),
    .B(_0840_),
    .C(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3918_ (.I(_0910_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3919_ (.I(_0943_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3920_ (.A1(_0854_),
    .A2(_0873_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3921_ (.A1(_0854_),
    .A2(_0868_),
    .A3(_0872_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3922_ (.A1(_0948_),
    .A2(_0832_),
    .B(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3923_ (.I(_0941_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3924_ (.A1(_0951_),
    .A2(_0937_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3925_ (.A1(_0947_),
    .A2(_0950_),
    .B(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3926_ (.I(_0890_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3927_ (.A1(_0954_),
    .A2(_0901_),
    .A3(_0904_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3928_ (.A1(_0946_),
    .A2(_0953_),
    .B(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3929_ (.I(\mod.pc_2[13] ),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_0780_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_0576_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3932_ (.I(_0572_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3933_ (.A1(\mod.registers.r13[13] ),
    .A2(_0959_),
    .B1(_0960_),
    .B2(\mod.registers.r6[13] ),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3934_ (.I(_0467_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_3171_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3936_ (.A1(\mod.registers.r7[13] ),
    .A2(_0962_),
    .B1(_0963_),
    .B2(\mod.registers.r3[13] ),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3937_ (.I(_0509_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3938_ (.A1(\mod.registers.r1[13] ),
    .A2(_0965_),
    .B(_0436_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_0460_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_0578_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3941_ (.A1(\mod.registers.r5[13] ),
    .A2(_0967_),
    .B1(_0968_),
    .B2(\mod.registers.r10[13] ),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3942_ (.A1(_0961_),
    .A2(_0964_),
    .A3(_0966_),
    .A4(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3943_ (.I(_0581_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3944_ (.I(_0571_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3945_ (.A1(\mod.registers.r8[13] ),
    .A2(_0971_),
    .B1(_0972_),
    .B2(\mod.registers.r2[13] ),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3946_ (.I(_0628_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3947_ (.I(_0626_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3948_ (.A1(\mod.registers.r4[13] ),
    .A2(_0974_),
    .B1(_0975_),
    .B2(\mod.registers.r11[13] ),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_0639_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_0516_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3951_ (.A1(\mod.registers.r9[13] ),
    .A2(_0977_),
    .B1(_0978_),
    .B2(\mod.registers.r12[13] ),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3952_ (.I(_0624_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3953_ (.I(_0518_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3954_ (.A1(\mod.registers.r14[13] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\mod.registers.r15[13] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3955_ (.A1(_0973_),
    .A2(_0976_),
    .A3(_0979_),
    .A4(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3956_ (.A1(_0970_),
    .A2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3957_ (.A1(_0957_),
    .A2(_0958_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3958_ (.I(_0804_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3959_ (.I(_0494_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3960_ (.I(_0548_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3961_ (.A1(\mod.registers.r7[13] ),
    .A2(_0987_),
    .B1(_0988_),
    .B2(\mod.registers.r11[13] ),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3962_ (.A1(\mod.registers.r12[13] ),
    .A2(_0893_),
    .B1(_0823_),
    .B2(\mod.registers.r2[13] ),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3963_ (.I(_0493_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3964_ (.I(_0480_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3965_ (.A1(\mod.registers.r10[13] ),
    .A2(_0991_),
    .B1(_0992_),
    .B2(\mod.registers.r13[13] ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3966_ (.A1(\mod.registers.r9[13] ),
    .A2(_0855_),
    .B1(_0863_),
    .B2(\mod.registers.r1[13] ),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3967_ (.A1(_0989_),
    .A2(_0990_),
    .A3(_0993_),
    .A4(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3968_ (.A1(\mod.registers.r5[13] ),
    .A2(_0559_),
    .B1(_0816_),
    .B2(\mod.registers.r6[13] ),
    .C1(\mod.registers.r14[13] ),
    .C2(_0820_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3969_ (.I(_0806_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3970_ (.A1(\mod.registers.r8[13] ),
    .A2(_0813_),
    .B1(_0997_),
    .B2(\mod.registers.r4[13] ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3971_ (.A1(\mod.registers.r15[13] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(\mod.registers.r3[13] ),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3972_ (.A1(_0996_),
    .A2(_0998_),
    .A3(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3973_ (.A1(_0995_),
    .A2(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3974_ (.A1(_0986_),
    .A2(_1001_),
    .B(_0827_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3975_ (.I(_0932_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3976_ (.A1(_0427_),
    .A2(_0829_),
    .B(_0902_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3977_ (.A1(_1003_),
    .A2(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3978_ (.A1(_1002_),
    .A2(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(_0985_),
    .A2(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3980_ (.A1(\mod.pc_2[13] ),
    .A2(_3127_),
    .B1(_0970_),
    .B2(_0983_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3981_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3982_ (.A1(_1009_),
    .A2(_1002_),
    .A3(_1005_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3983_ (.A1(_1007_),
    .A2(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3984_ (.A1(\mod.pc_2[12] ),
    .A2(_0834_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3985_ (.A1(\mod.registers.r11[12] ),
    .A2(_0975_),
    .B1(_0963_),
    .B2(\mod.registers.r3[12] ),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3986_ (.A1(\mod.registers.r6[12] ),
    .A2(_0960_),
    .B1(_0968_),
    .B2(\mod.registers.r10[12] ),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3987_ (.A1(\mod.registers.r9[12] ),
    .A2(_0977_),
    .B(_0522_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3988_ (.A1(\mod.registers.r4[12] ),
    .A2(_0974_),
    .B1(_0980_),
    .B2(\mod.registers.r14[12] ),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3989_ (.A1(_1013_),
    .A2(_1014_),
    .A3(_1015_),
    .A4(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3990_ (.A1(\mod.registers.r15[12] ),
    .A2(_0981_),
    .B1(_0978_),
    .B2(\mod.registers.r12[12] ),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3991_ (.A1(\mod.registers.r13[12] ),
    .A2(_0959_),
    .B1(_0965_),
    .B2(\mod.registers.r1[12] ),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3992_ (.A1(\mod.registers.r8[12] ),
    .A2(_0971_),
    .B1(_0962_),
    .B2(\mod.registers.r7[12] ),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3993_ (.A1(\mod.registers.r5[12] ),
    .A2(_0967_),
    .B1(_0972_),
    .B2(\mod.registers.r2[12] ),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3994_ (.A1(_1018_),
    .A2(_1019_),
    .A3(_1020_),
    .A4(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3995_ (.A1(_1017_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3996_ (.A1(_1012_),
    .A2(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3997_ (.A1(\mod.registers.r10[12] ),
    .A2(_0991_),
    .B1(_0997_),
    .B2(\mod.registers.r4[12] ),
    .C1(_0988_),
    .C2(\mod.registers.r11[12] ),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3998_ (.A1(\mod.registers.r9[12] ),
    .A2(_0805_),
    .B1(_0987_),
    .B2(\mod.registers.r7[12] ),
    .C1(_0821_),
    .C2(\mod.registers.r14[12] ),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3999_ (.A1(\mod.registers.r1[12] ),
    .A2(_0824_),
    .B1(_0992_),
    .B2(\mod.registers.r13[12] ),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4000_ (.A1(\mod.registers.r5[12] ),
    .A2(_0819_),
    .B1(_0858_),
    .B2(\mod.registers.r8[12] ),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4001_ (.A1(\mod.registers.r15[12] ),
    .A2(_0558_),
    .B1(_0898_),
    .B2(\mod.registers.r6[12] ),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4002_ (.A1(\mod.registers.r12[12] ),
    .A2(_0555_),
    .B1(_0865_),
    .B2(\mod.registers.r2[12] ),
    .C1(_0859_),
    .C2(\mod.registers.r3[12] ),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4003_ (.A1(_1028_),
    .A2(_1029_),
    .A3(_1030_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4004_ (.A1(_1025_),
    .A2(_1026_),
    .A3(_1027_),
    .A4(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4005_ (.A1(_0986_),
    .A2(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4006_ (.I(_0829_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4007_ (.I(_0902_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4008_ (.A1(_0524_),
    .A2(_1034_),
    .B(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4009_ (.I(_0456_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4010_ (.A1(_0827_),
    .A2(_1033_),
    .B1(_1036_),
    .B2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4011_ (.A1(_1024_),
    .A2(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4012_ (.A1(_1024_),
    .A2(_1038_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4013_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4014_ (.A1(_0945_),
    .A2(_0956_),
    .B(_1011_),
    .C(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4015_ (.A1(_1009_),
    .A2(_1006_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4016_ (.I(\mod.pc_2[12] ),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4017_ (.A1(_1044_),
    .A2(_0958_),
    .B(_1023_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4018_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4019_ (.A1(_1011_),
    .A2(_1046_),
    .A3(_1038_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4020_ (.A1(_1043_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4021_ (.A1(\mod.registers.r7[14] ),
    .A2(_0962_),
    .B1(_0960_),
    .B2(\mod.registers.r6[14] ),
    .C1(_0959_),
    .C2(\mod.registers.r13[14] ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4022_ (.A1(\mod.registers.r14[14] ),
    .A2(_0980_),
    .B1(_0965_),
    .B2(\mod.registers.r1[14] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4023_ (.A1(\mod.registers.r4[14] ),
    .A2(_0974_),
    .B1(_0975_),
    .B2(\mod.registers.r11[14] ),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4024_ (.A1(_1049_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4025_ (.A1(\mod.registers.r9[14] ),
    .A2(_0977_),
    .B1(_0967_),
    .B2(\mod.registers.r5[14] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4026_ (.A1(\mod.registers.r15[14] ),
    .A2(_0981_),
    .B1(_0978_),
    .B2(\mod.registers.r12[14] ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4027_ (.A1(\mod.registers.r8[14] ),
    .A2(_0971_),
    .B1(_0968_),
    .B2(\mod.registers.r10[14] ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4028_ (.A1(\mod.registers.r3[14] ),
    .A2(_0963_),
    .B1(_0972_),
    .B2(\mod.registers.r2[14] ),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4029_ (.A1(_1053_),
    .A2(_1054_),
    .A3(_1055_),
    .A4(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4030_ (.A1(_1052_),
    .A2(_1057_),
    .B(_0834_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4031_ (.I(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4032_ (.A1(\mod.registers.r13[14] ),
    .A2(_0992_),
    .B1(_0997_),
    .B2(\mod.registers.r4[14] ),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4033_ (.A1(\mod.registers.r9[14] ),
    .A2(_0805_),
    .B1(_0987_),
    .B2(\mod.registers.r7[14] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4034_ (.A1(\mod.registers.r5[14] ),
    .A2(_0819_),
    .B1(_0823_),
    .B2(\mod.registers.r2[14] ),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4035_ (.A1(\mod.registers.r10[14] ),
    .A2(_0991_),
    .B1(_0824_),
    .B2(\mod.registers.r1[14] ),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4036_ (.A1(_1060_),
    .A2(_1061_),
    .A3(_1062_),
    .A4(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4037_ (.A1(\mod.registers.r8[14] ),
    .A2(_0813_),
    .B1(_0898_),
    .B2(\mod.registers.r6[14] ),
    .C1(_0893_),
    .C2(\mod.registers.r12[14] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4038_ (.A1(\mod.registers.r14[14] ),
    .A2(_0821_),
    .B1(_0988_),
    .B2(\mod.registers.r11[14] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4039_ (.A1(\mod.registers.r15[14] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(\mod.registers.r3[14] ),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4040_ (.A1(_1065_),
    .A2(_1066_),
    .A3(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4041_ (.A1(_1064_),
    .A2(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4042_ (.A1(_0986_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4043_ (.A1(_3196_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4044_ (.I(_3106_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4045_ (.A1(_0441_),
    .A2(_1072_),
    .A3(_3165_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4046_ (.I(_3194_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4047_ (.A1(_1074_),
    .A2(_0986_),
    .B(_1070_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4048_ (.A1(_1059_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4049_ (.A1(_1059_),
    .A2(_1071_),
    .A3(_1073_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4050_ (.I(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4051_ (.A1(_1042_),
    .A2(_1048_),
    .B(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4052_ (.I(_1058_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4053_ (.A1(_1080_),
    .A2(_1075_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4054_ (.I(_1003_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4055_ (.A1(\mod.registers.r1[15] ),
    .A2(_0965_),
    .B1(_0963_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4056_ (.A1(\mod.registers.r7[15] ),
    .A2(_0962_),
    .B1(_0967_),
    .B2(\mod.registers.r5[15] ),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4057_ (.A1(_1083_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4058_ (.A1(\mod.registers.r6[15] ),
    .A2(_0960_),
    .B1(_0978_),
    .B2(\mod.registers.r12[15] ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4059_ (.A1(\mod.registers.r9[15] ),
    .A2(_0977_),
    .B1(_0968_),
    .B2(\mod.registers.r10[15] ),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4060_ (.A1(\mod.registers.r13[15] ),
    .A2(_0959_),
    .B1(_0980_),
    .B2(\mod.registers.r14[15] ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4061_ (.A1(\mod.registers.r4[15] ),
    .A2(_0974_),
    .B1(_0972_),
    .B2(\mod.registers.r2[15] ),
    .C1(_0975_),
    .C2(\mod.registers.r11[15] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4062_ (.A1(\mod.registers.r8[15] ),
    .A2(_0971_),
    .B1(_0981_),
    .B2(\mod.registers.r15[15] ),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4063_ (.A1(_1088_),
    .A2(_1089_),
    .A3(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4064_ (.A1(_1085_),
    .A2(_1086_),
    .A3(_1087_),
    .A4(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4065_ (.A1(_1082_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4066_ (.I(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4067_ (.A1(\mod.registers.r10[15] ),
    .A2(_0991_),
    .B1(_0824_),
    .B2(\mod.registers.r1[15] ),
    .C1(_0997_),
    .C2(\mod.registers.r4[15] ),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4068_ (.A1(\mod.registers.r13[15] ),
    .A2(_0992_),
    .B1(_0987_),
    .B2(\mod.registers.r7[15] ),
    .C1(_0821_),
    .C2(\mod.registers.r14[15] ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4069_ (.A1(\mod.registers.r9[15] ),
    .A2(_0805_),
    .B1(_0988_),
    .B2(\mod.registers.r11[15] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4070_ (.A1(_1095_),
    .A2(_1096_),
    .A3(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4071_ (.A1(\mod.registers.r5[15] ),
    .A2(_0819_),
    .B1(_0813_),
    .B2(\mod.registers.r8[15] ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4072_ (.A1(\mod.registers.r15[15] ),
    .A2(_0810_),
    .B1(_0898_),
    .B2(\mod.registers.r6[15] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4073_ (.A1(\mod.registers.r2[15] ),
    .A2(_0823_),
    .B1(_0811_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4074_ (.A1(_1099_),
    .A2(_1100_),
    .A3(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4075_ (.A1(\mod.registers.r12[15] ),
    .A2(_0893_),
    .B(_1098_),
    .C(_1102_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4076_ (.A1(_0539_),
    .A2(_1103_),
    .B(_3196_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4077_ (.I(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4078_ (.A1(_0413_),
    .A2(_1034_),
    .B(_1035_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4079_ (.A1(_1082_),
    .A2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4080_ (.A1(_1094_),
    .A2(_1105_),
    .A3(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4081_ (.A1(_1085_),
    .A2(_1086_),
    .A3(_1087_),
    .A4(_1091_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4082_ (.I(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4083_ (.A1(_1110_),
    .A2(_1104_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4084_ (.A1(_1108_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4085_ (.I(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4086_ (.A1(_1079_),
    .A2(_1081_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4087_ (.A1(_1113_),
    .A2(_1079_),
    .A3(_1081_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4088_ (.A1(\mod.funct7[1] ),
    .A2(_3114_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4089_ (.A1(_3120_),
    .A2(_3109_),
    .B(_1116_),
    .C(_3111_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4090_ (.A1(_3117_),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4091_ (.I(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4092_ (.I(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4093_ (.I(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4094_ (.A1(_1114_),
    .A2(_1115_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4095_ (.A1(_3117_),
    .A2(_1117_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4096_ (.I(_1123_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4097_ (.I(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4098_ (.I(_1039_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4099_ (.I(_1010_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4100_ (.A1(_1007_),
    .A2(_1126_),
    .B(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_0598_),
    .A2(_0602_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4102_ (.A1(_0703_),
    .A2(_0705_),
    .A3(_0725_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4103_ (.I(_0747_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4104_ (.I(_0748_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4105_ (.I(\mod.pc_2[0] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4106_ (.A1(_0749_),
    .A2(_0750_),
    .A3(_0751_),
    .A4(_0752_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4107_ (.A1(_0754_),
    .A2(_0755_),
    .A3(_0757_),
    .A4(_0758_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4108_ (.A1(_1133_),
    .A2(_0932_),
    .B1(_1134_),
    .B2(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4109_ (.A1(_1131_),
    .A2(_1132_),
    .A3(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4110_ (.A1(_1130_),
    .A2(_1137_),
    .B(_0735_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4111_ (.I(_0674_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4112_ (.I(_0681_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4113_ (.A1(_0770_),
    .A2(_0771_),
    .A3(_1139_),
    .A4(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4114_ (.A1(_0619_),
    .A2(_0620_),
    .A3(_0642_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4115_ (.A1(_1142_),
    .A2(_1140_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4116_ (.A1(_1138_),
    .A2(_1141_),
    .B(_1143_),
    .C(_1139_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4117_ (.A1(_0593_),
    .A2(_0543_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4118_ (.A1(_1145_),
    .A2(_0777_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4119_ (.I(_0598_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4120_ (.I(_0602_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4121_ (.I(_0521_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4122_ (.I(_0543_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4123_ (.A1(_1149_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4124_ (.A1(_1149_),
    .A2(_1150_),
    .B(_0776_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4125_ (.A1(_1147_),
    .A2(_1148_),
    .A3(_1151_),
    .A4(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4126_ (.A1(_1129_),
    .A2(_1144_),
    .A3(_1146_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4127_ (.I(_0597_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4128_ (.A1(_1155_),
    .A2(_0450_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(_0600_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4130_ (.A1(_1155_),
    .A2(_0450_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4131_ (.A1(_1156_),
    .A2(_1157_),
    .B(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4132_ (.A1(_0832_),
    .A2(_0839_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4133_ (.A1(_0877_),
    .A2(_0910_),
    .A3(_0947_),
    .A4(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_1154_),
    .A2(_1159_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4135_ (.I(_0922_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4136_ (.A1(_1163_),
    .A2(_0937_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4137_ (.I(_0854_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4138_ (.A1(_1165_),
    .A2(_0873_),
    .B(_0803_),
    .C(_0838_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4139_ (.A1(_0874_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4140_ (.A1(_1164_),
    .A2(_1167_),
    .B(_0906_),
    .C(_0938_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_0909_),
    .A2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4142_ (.A1(_1162_),
    .A2(_1169_),
    .B(_1011_),
    .C(_1041_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4143_ (.A1(_1128_),
    .A2(_1170_),
    .B(_1078_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4144_ (.A1(_1076_),
    .A2(_1171_),
    .B(_1112_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4145_ (.A1(_1112_),
    .A2(_1076_),
    .A3(_1171_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4146_ (.A1(_1125_),
    .A2(_1172_),
    .A3(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4147_ (.I(\mod.funct3[1] ),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4148_ (.A1(_1175_),
    .A2(_3122_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4149_ (.I(\mod.funct3[2] ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4150_ (.A1(_0437_),
    .A2(_0569_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4151_ (.A1(_1177_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4152_ (.I(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4153_ (.A1(_1176_),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4154_ (.I(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4155_ (.A1(_1003_),
    .A2(_0660_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4156_ (.I(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4157_ (.I(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4158_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4159_ (.A1(_0932_),
    .A2(_0729_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4160_ (.I(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4161_ (.A1(_0780_),
    .A2(_0765_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4162_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4163_ (.A1(_1188_),
    .A2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4164_ (.I(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4165_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_0645_),
    .A2(_0525_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4167_ (.A1(_0562_),
    .A2(_0738_),
    .A3(_0746_),
    .B(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4168_ (.I(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4169_ (.A1(_0834_),
    .A2(_1109_),
    .A3(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4170_ (.A1(_1193_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4171_ (.A1(_1092_),
    .A2(_1118_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4172_ (.I(_0567_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4173_ (.I(_0683_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4174_ (.A1(_1200_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_1199_),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4176_ (.I(_0706_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4177_ (.I(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4178_ (.A1(_0569_),
    .A2(_1195_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4179_ (.I(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4181_ (.I(_1190_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4182_ (.A1(_1208_),
    .A2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(_1205_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4184_ (.A1(_1211_),
    .A2(_1199_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4185_ (.A1(_1186_),
    .A2(_1198_),
    .B(_1203_),
    .C(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4186_ (.A1(_1182_),
    .A2(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4187_ (.I(_1175_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4188_ (.I(_3122_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4189_ (.A1(_1215_),
    .A2(_1216_),
    .A3(_1179_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4190_ (.I(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4191_ (.A1(_3120_),
    .A2(_3128_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4192_ (.I(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4193_ (.A1(\mod.funct3[1] ),
    .A2(_3122_),
    .A3(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4194_ (.I(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4195_ (.I(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4196_ (.A1(_1111_),
    .A2(_1223_),
    .B(_3131_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_1220_),
    .A2(_3123_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4198_ (.A1(_1112_),
    .A2(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4199_ (.A1(_1108_),
    .A2(_1218_),
    .B(_1224_),
    .C(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4200_ (.I(_1184_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4201_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4202_ (.I(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4203_ (.I(_1196_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4204_ (.A1(_1037_),
    .A2(_1058_),
    .A3(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4205_ (.A1(_1197_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4206_ (.I(_0706_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4207_ (.I(_1189_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4208_ (.A1(_1234_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4209_ (.I(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4210_ (.I(_1206_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4211_ (.I(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4212_ (.A1(_1131_),
    .A2(_1132_),
    .B(_1008_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4213_ (.A1(_1239_),
    .A2(_1046_),
    .B(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4214_ (.I(_0621_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4215_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4216_ (.I(_1188_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_1238_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4218_ (.I(_0908_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4219_ (.A1(_1246_),
    .A2(_1208_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4220_ (.A1(_1163_),
    .A2(_1245_),
    .B(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4221_ (.I(_0803_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4222_ (.A1(_1131_),
    .A2(_1132_),
    .A3(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4223_ (.A1(_0875_),
    .A2(_1245_),
    .B(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4224_ (.A1(_1244_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4225_ (.A1(_1244_),
    .A2(_1248_),
    .B(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4226_ (.A1(_1243_),
    .A2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4227_ (.A1(_1193_),
    .A2(_1233_),
    .B1(_1237_),
    .B2(_1241_),
    .C(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4228_ (.I(_1201_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4229_ (.I(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4230_ (.A1(_1003_),
    .A2(_1196_),
    .A3(_1136_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4231_ (.I(_1131_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4232_ (.I(_1132_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4233_ (.A1(_1259_),
    .A2(_1260_),
    .B(_0726_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4234_ (.A1(_1258_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4235_ (.I(_0673_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4236_ (.A1(_0747_),
    .A2(_0748_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4237_ (.I(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4238_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4239_ (.A1(_1037_),
    .A2(_1196_),
    .A3(_0643_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4240_ (.A1(_1263_),
    .A2(_1266_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4241_ (.I(_0706_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4242_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4243_ (.I0(_1262_),
    .I1(_1268_),
    .S(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4244_ (.I(_0593_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4245_ (.I(_0589_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4246_ (.I0(_1272_),
    .I1(_1273_),
    .S(_1238_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4247_ (.A1(_1082_),
    .A2(_1231_),
    .B(_0597_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4248_ (.A1(_0599_),
    .A2(_1266_),
    .B(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4249_ (.I0(_1274_),
    .I1(_1276_),
    .S(_1270_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4250_ (.I(_0621_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4251_ (.I0(_1271_),
    .I1(_1277_),
    .S(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4252_ (.A1(_1257_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4253_ (.A1(_1177_),
    .A2(_3129_),
    .A3(_1176_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4254_ (.A1(_1230_),
    .A2(_1255_),
    .B(_1280_),
    .C(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4255_ (.A1(_1214_),
    .A2(_1227_),
    .A3(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4256_ (.A1(_1177_),
    .A2(_3129_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4257_ (.A1(_3118_),
    .A2(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4258_ (.I(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4259_ (.A1(_1114_),
    .A2(_1115_),
    .B(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4260_ (.A1(_3132_),
    .A2(_1122_),
    .A3(_1174_),
    .B1(_1283_),
    .B2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4261_ (.I(_1124_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4262_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4263_ (.I(_0938_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4264_ (.I(_0832_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4265_ (.I(_0840_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4266_ (.A1(_0605_),
    .A2(_0778_),
    .B(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4267_ (.A1(_1292_),
    .A2(_1294_),
    .B(_0877_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4268_ (.A1(_1291_),
    .A2(_0942_),
    .B1(_0949_),
    .B2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4269_ (.I(_0946_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4270_ (.A1(_0952_),
    .A2(_1296_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4271_ (.A1(_1297_),
    .A2(_0952_),
    .A3(_1296_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4272_ (.A1(_1290_),
    .A2(_1298_),
    .A3(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4273_ (.I(_1120_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4274_ (.I(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4275_ (.I(_0948_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4276_ (.A1(_1154_),
    .A2(_1159_),
    .B(_1303_),
    .C(_1293_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4277_ (.A1(_1167_),
    .A2(_1304_),
    .B(_0947_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4278_ (.A1(_1163_),
    .A2(_0937_),
    .B(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4279_ (.A1(_1297_),
    .A2(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4280_ (.A1(_1302_),
    .A2(_1307_),
    .B(_3132_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4281_ (.I(_1286_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4282_ (.A1(_1298_),
    .A2(_1299_),
    .B(_1309_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4283_ (.I(\mod.funct3[0] ),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4284_ (.A1(_1215_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4285_ (.A1(_1180_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4286_ (.I(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4288_ (.A1(_0954_),
    .A2(_0905_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4289_ (.I(_1311_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4290_ (.A1(_3118_),
    .A2(_1317_),
    .A3(_1219_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4291_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4292_ (.I(_1222_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4293_ (.A1(_1316_),
    .A2(_1319_),
    .B1(_1320_),
    .B2(_0906_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4294_ (.I(_1229_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4295_ (.I(_1242_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(_1323_),
    .A2(_1271_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4297_ (.I(_1323_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(_1209_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4299_ (.A1(_1326_),
    .A2(_1277_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4300_ (.A1(_1325_),
    .A2(_1253_),
    .B(_1327_),
    .C(_1186_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4301_ (.I(_1215_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4302_ (.A1(_1329_),
    .A2(_1216_),
    .A3(_1284_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4303_ (.I(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4304_ (.A1(_1322_),
    .A2(_1324_),
    .B(_1328_),
    .C(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4305_ (.A1(_1297_),
    .A2(_1315_),
    .B(_1321_),
    .C(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4306_ (.I(_1182_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4307_ (.I(_1264_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4308_ (.I0(_1080_),
    .I1(_1009_),
    .I2(_1024_),
    .I3(_1246_),
    .S0(_1335_),
    .S1(_1234_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4309_ (.I(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4310_ (.I(_1187_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4311_ (.I(_1338_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4312_ (.A1(_1339_),
    .A2(_1242_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4313_ (.A1(_1323_),
    .A2(_1337_),
    .B1(_1340_),
    .B2(_1197_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_1326_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4315_ (.A1(_1244_),
    .A2(_1239_),
    .B(_1342_),
    .C(_1199_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(_1203_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4317_ (.A1(_1322_),
    .A2(_1341_),
    .B(_1343_),
    .C(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_1334_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4319_ (.A1(_1333_),
    .A2(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4320_ (.A1(_1300_),
    .A2(_1308_),
    .B(_1310_),
    .C(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4321_ (.A1(_1119_),
    .A2(_3130_),
    .B(_1285_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4322_ (.A1(_1007_),
    .A2(_1010_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4323_ (.I(_1041_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4324_ (.A1(_0945_),
    .A2(_0956_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4325_ (.A1(_1046_),
    .A2(_1038_),
    .B1(_1351_),
    .B2(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4326_ (.A1(_1350_),
    .A2(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4327_ (.I(_1338_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4328_ (.A1(_1355_),
    .A2(_1197_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4329_ (.A1(_1232_),
    .A2(_1240_),
    .B(_1269_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4330_ (.I(_1190_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4331_ (.A1(_1356_),
    .A2(_1357_),
    .B(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4332_ (.A1(_0729_),
    .A2(_0765_),
    .B(_0958_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(_1360_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_1093_),
    .A2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4335_ (.A1(_1200_),
    .A2(_1289_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4336_ (.A1(_1210_),
    .A2(_1362_),
    .A3(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4337_ (.A1(_1359_),
    .A2(_1364_),
    .B(_1257_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4338_ (.A1(_1344_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4339_ (.I(_1256_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4340_ (.I(_1264_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4341_ (.A1(_1263_),
    .A2(_1368_),
    .B(_1267_),
    .C(_1234_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4342_ (.A1(_1270_),
    .A2(_1274_),
    .B(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4343_ (.I(_1204_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(_1371_),
    .A2(_1262_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4345_ (.I(_1189_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4346_ (.I0(_1370_),
    .I1(_1372_),
    .S(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4347_ (.A1(_1367_),
    .A2(_1331_),
    .A3(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4348_ (.A1(_1010_),
    .A2(_1218_),
    .B1(_1314_),
    .B2(_1350_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4349_ (.I(_1242_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4350_ (.I0(_1276_),
    .I1(_1251_),
    .S(_1371_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4351_ (.A1(_1201_),
    .A2(_1281_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4352_ (.I(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4353_ (.A1(_1248_),
    .A2(_1237_),
    .B1(_1241_),
    .B2(_1192_),
    .C(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4354_ (.A1(_1377_),
    .A2(_1378_),
    .B(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4355_ (.A1(_1007_),
    .A2(_1223_),
    .B(_1376_),
    .C(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4356_ (.A1(_1182_),
    .A2(_1366_),
    .B(_1375_),
    .C(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4357_ (.I(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4358_ (.I(_1126_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4359_ (.A1(_1162_),
    .A2(_1169_),
    .B(_1351_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4360_ (.A1(_1350_),
    .A2(_1386_),
    .A3(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4361_ (.A1(_1124_),
    .A2(_3130_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4362_ (.A1(_1386_),
    .A2(_1387_),
    .B(_1350_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4363_ (.A1(_1388_),
    .A2(_1389_),
    .A3(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4364_ (.A1(_1349_),
    .A2(_1354_),
    .B(_1385_),
    .C(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4365_ (.A1(_0877_),
    .A2(_1292_),
    .A3(_1294_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4366_ (.A1(_1295_),
    .A2(_1393_),
    .B(_1121_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4367_ (.A1(_1249_),
    .A2(_0838_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4368_ (.A1(_1154_),
    .A2(_1159_),
    .B(_1293_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4369_ (.A1(_1395_),
    .A2(_1396_),
    .B(_1303_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4370_ (.A1(_1303_),
    .A2(_1395_),
    .A3(_1396_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4371_ (.I(_1177_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4372_ (.A1(_1399_),
    .A2(_1312_),
    .B(_1178_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4373_ (.I(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4374_ (.I(_1401_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4375_ (.A1(_1125_),
    .A2(_1397_),
    .A3(_1398_),
    .B(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4376_ (.A1(_1399_),
    .A2(_1215_),
    .A3(_3129_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4377_ (.I(_1404_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4378_ (.A1(_1405_),
    .A2(_1295_),
    .A3(_1393_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4379_ (.I(_1235_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4380_ (.I(_1407_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4381_ (.I0(_1165_),
    .I1(_0954_),
    .I2(_0922_),
    .I3(_1045_),
    .S0(_1338_),
    .S1(_1207_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4382_ (.A1(_1356_),
    .A2(_1357_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4383_ (.A1(_1326_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4384_ (.I(_1201_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4385_ (.A1(_1408_),
    .A2(_1409_),
    .B(_1411_),
    .C(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4386_ (.I(_1335_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4387_ (.A1(_1109_),
    .A2(_1355_),
    .A3(_1235_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4388_ (.A1(_1414_),
    .A2(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4389_ (.A1(_1119_),
    .A2(_1202_),
    .A3(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4390_ (.A1(_1344_),
    .A2(_1413_),
    .A3(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_1262_),
    .A2(_1192_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4392_ (.A1(_1243_),
    .A2(_1370_),
    .B(_1256_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4393_ (.A1(_1377_),
    .A2(_1378_),
    .B(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4394_ (.A1(_1186_),
    .A2(_1419_),
    .B(_1421_),
    .C(_1330_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4395_ (.A1(_1303_),
    .A2(_1314_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(_0876_),
    .A2(_1217_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4397_ (.A1(_0874_),
    .A2(_1223_),
    .B(_1423_),
    .C(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4398_ (.A1(_1182_),
    .A2(_1418_),
    .B(_1422_),
    .C(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4399_ (.A1(_1394_),
    .A2(_1403_),
    .B(_1406_),
    .C(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4400_ (.I(_1148_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4401_ (.A1(_1190_),
    .A2(_0769_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4402_ (.A1(_1139_),
    .A2(_1140_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4403_ (.A1(_1184_),
    .A2(_1263_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4404_ (.A1(_1429_),
    .A2(_1430_),
    .B(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4405_ (.A1(_1188_),
    .A2(_0733_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4406_ (.A1(_0958_),
    .A2(_0729_),
    .B(_0733_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4407_ (.A1(_1130_),
    .A2(_1434_),
    .B(_1258_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4408_ (.A1(_0770_),
    .A2(_0771_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4409_ (.A1(_1433_),
    .A2(_1435_),
    .B(_1436_),
    .C(_1430_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4410_ (.A1(_0567_),
    .A2(_0588_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_0589_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4412_ (.A1(_0775_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4413_ (.A1(_1438_),
    .A2(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4414_ (.A1(_1432_),
    .A2(_1437_),
    .B(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4415_ (.A1(_1200_),
    .A2(_1273_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4416_ (.A1(_1442_),
    .A2(_1443_),
    .B(_1145_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(_0594_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4418_ (.A1(_1428_),
    .A2(_1445_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4419_ (.I(_1144_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4420_ (.A1(_1151_),
    .A2(_1152_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4421_ (.A1(_1447_),
    .A2(_1146_),
    .B(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4422_ (.A1(_1428_),
    .A2(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4423_ (.A1(_1125_),
    .A2(_1450_),
    .B(_1402_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4424_ (.A1(_1290_),
    .A2(_1446_),
    .B(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4425_ (.A1(_1109_),
    .A2(_0775_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4426_ (.I(_1183_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4427_ (.A1(_1093_),
    .A2(_1200_),
    .A3(_1454_),
    .A4(_1361_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4428_ (.A1(_0775_),
    .A2(_1184_),
    .B(_1123_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4429_ (.A1(_1453_),
    .A2(_1455_),
    .B(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4430_ (.I0(_0954_),
    .I1(_1163_),
    .I2(_0985_),
    .I3(_1045_),
    .S0(_1368_),
    .S1(_1355_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4431_ (.A1(_1377_),
    .A2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4432_ (.I(_0473_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4433_ (.I0(_1165_),
    .I1(_1155_),
    .I2(_1249_),
    .I3(_1460_),
    .S0(_1269_),
    .S1(_1266_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4434_ (.A1(_1408_),
    .A2(_1461_),
    .B(_1257_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4435_ (.A1(_1110_),
    .A2(_1414_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4436_ (.A1(_1080_),
    .A2(_1414_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_1192_),
    .A2(_1464_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4438_ (.A1(_1459_),
    .A2(_1462_),
    .B1(_1465_),
    .B2(_1257_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4439_ (.A1(_1457_),
    .A2(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4440_ (.I(_1216_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4441_ (.A1(_1329_),
    .A2(_1468_),
    .A3(_1220_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4442_ (.A1(_1329_),
    .A2(_0600_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4443_ (.A1(_1468_),
    .A2(_1157_),
    .B(_0601_),
    .C(_1180_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4444_ (.A1(_1263_),
    .A2(_1259_),
    .A3(_1260_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4445_ (.A1(_1273_),
    .A2(_1245_),
    .B(_1472_),
    .C(_1244_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4446_ (.A1(_1149_),
    .A2(_1259_),
    .A3(_1260_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4447_ (.A1(_1460_),
    .A2(_1245_),
    .B(_1474_),
    .C(_1371_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4448_ (.A1(_1473_),
    .A2(_1475_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4449_ (.A1(_1037_),
    .A2(_0726_),
    .A3(_1231_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4450_ (.A1(_1368_),
    .A2(_0769_),
    .B(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4451_ (.A1(_1238_),
    .A2(_0760_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4452_ (.I0(_1478_),
    .I1(_1479_),
    .S(_1339_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(_1408_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4454_ (.A1(_1408_),
    .A2(_1476_),
    .B(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4455_ (.A1(_1454_),
    .A2(_1330_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4456_ (.A1(_1470_),
    .A2(_1471_),
    .B1(_1482_),
    .B2(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4457_ (.A1(_1286_),
    .A2(_1446_),
    .B1(_1467_),
    .B2(_1469_),
    .C(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4458_ (.A1(_0840_),
    .A2(_1154_),
    .A3(_1159_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4459_ (.A1(_1396_),
    .A2(_1486_),
    .B(_1289_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4460_ (.A1(_0605_),
    .A2(_0778_),
    .B(_1160_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4461_ (.A1(_1272_),
    .A2(_1150_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4462_ (.A1(_1145_),
    .A2(_1443_),
    .B(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4463_ (.A1(_0451_),
    .A2(_0505_),
    .B(_0604_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4464_ (.A1(_1147_),
    .A2(_1148_),
    .A3(_1490_),
    .B(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(_0544_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4466_ (.A1(_1147_),
    .A2(_1148_),
    .A3(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4467_ (.A1(_1432_),
    .A2(_1437_),
    .B(_1494_),
    .C(_1441_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4468_ (.A1(_1492_),
    .A2(_1495_),
    .A3(_1293_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4469_ (.A1(_1120_),
    .A2(_1488_),
    .A3(_1496_),
    .B(_1401_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4470_ (.A1(_1488_),
    .A2(_1496_),
    .B(_1404_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4471_ (.A1(_1329_),
    .A2(_1395_),
    .B1(_1160_),
    .B2(_1468_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4472_ (.I0(_1092_),
    .I1(_1058_),
    .I2(_1009_),
    .I3(_1024_),
    .S0(_1264_),
    .S1(_1204_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4473_ (.I0(_0875_),
    .I1(_1246_),
    .I2(_0837_),
    .I3(_0951_),
    .S0(_1338_),
    .S1(_1265_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4474_ (.I0(_1500_),
    .I1(_1501_),
    .S(_0621_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4475_ (.A1(_1229_),
    .A2(_1502_),
    .B(_1203_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4476_ (.I(_1181_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4477_ (.I0(_1439_),
    .I1(_0684_),
    .I2(_0643_),
    .I3(_0726_),
    .S0(_1206_),
    .S1(_1188_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_1407_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4479_ (.I0(_1460_),
    .I1(_1272_),
    .S(_1207_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4480_ (.I0(_1155_),
    .I1(_1249_),
    .S(_1265_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4481_ (.I0(_1507_),
    .I1(_1508_),
    .S(_1234_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4482_ (.A1(_1278_),
    .A2(_1509_),
    .B(_1228_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(_0683_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4484_ (.A1(_1082_),
    .A2(_1231_),
    .B(_1136_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4485_ (.A1(_1361_),
    .A2(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4486_ (.A1(_1511_),
    .A2(_1513_),
    .B(_1281_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4487_ (.A1(_1506_),
    .A2(_1510_),
    .B(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4488_ (.A1(_1220_),
    .A2(_1499_),
    .B1(_1503_),
    .B2(_1504_),
    .C(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4489_ (.A1(_1487_),
    .A2(_1497_),
    .B(_1498_),
    .C(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4490_ (.I(_0777_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4491_ (.A1(_0686_),
    .A2(_0773_),
    .B(_1518_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4492_ (.A1(_1493_),
    .A2(_1519_),
    .A3(_0590_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4493_ (.A1(_1444_),
    .A2(_1520_),
    .B(_1120_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4494_ (.A1(_1518_),
    .A2(_1447_),
    .B(_0776_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4495_ (.A1(_1493_),
    .A2(_1522_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4496_ (.A1(_1125_),
    .A2(_1523_),
    .B(_1401_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4497_ (.A1(_1405_),
    .A2(_1444_),
    .A3(_1520_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4498_ (.I0(_1460_),
    .I1(_1272_),
    .S(_1335_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4499_ (.A1(_1275_),
    .A2(_1250_),
    .B(_1371_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4500_ (.A1(_1205_),
    .A2(_1526_),
    .B(_1527_),
    .C(_1407_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4501_ (.A1(_1243_),
    .A2(_1409_),
    .B(_1256_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4502_ (.A1(_1210_),
    .A2(_1453_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4503_ (.A1(_1185_),
    .A2(_1359_),
    .B1(_1457_),
    .B2(_1530_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4504_ (.A1(_1528_),
    .A2(_1529_),
    .B(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4505_ (.A1(_1149_),
    .A2(_1150_),
    .A3(_1221_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4506_ (.A1(_1151_),
    .A2(_1217_),
    .B1(_1313_),
    .B2(_1493_),
    .C(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4507_ (.A1(_1380_),
    .A2(_1374_),
    .B(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4508_ (.A1(_1504_),
    .A2(_1532_),
    .B(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4509_ (.A1(_1521_),
    .A2(_1524_),
    .B(_1525_),
    .C(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_0761_),
    .A2(_1512_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4511_ (.I(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4512_ (.A1(_1511_),
    .A2(_1502_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4513_ (.I(_1453_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4514_ (.A1(_1119_),
    .A2(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4515_ (.I0(_0597_),
    .I1(_0473_),
    .I2(_0593_),
    .I3(_1439_),
    .S0(_1265_),
    .S1(_1204_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4516_ (.I0(_0684_),
    .I1(_0643_),
    .S(_1368_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4517_ (.A1(_1259_),
    .A2(_1260_),
    .B(_1136_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4518_ (.A1(_1360_),
    .A2(_1477_),
    .A3(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4519_ (.A1(_1358_),
    .A2(_1543_),
    .B1(_1544_),
    .B2(_1236_),
    .C(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(_1185_),
    .A2(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4521_ (.A1(_1540_),
    .A2(_1542_),
    .A3(_1548_),
    .B(_1181_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4522_ (.A1(_1404_),
    .A2(_1313_),
    .B(_1538_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4523_ (.A1(_1222_),
    .A2(_1137_),
    .B1(_1545_),
    .B2(_1319_),
    .C(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4524_ (.A1(_1483_),
    .A2(_1513_),
    .B(_1551_),
    .C(_1400_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4525_ (.A1(_1401_),
    .A2(_1539_),
    .B1(_1549_),
    .B2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4526_ (.A1(_1355_),
    .A2(_1275_),
    .A3(_1250_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4527_ (.A1(_1339_),
    .A2(_1526_),
    .B(_1554_),
    .C(_1209_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4528_ (.A1(_1261_),
    .A2(_1267_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4529_ (.I0(_1439_),
    .I1(_0684_),
    .S(_1335_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4530_ (.A1(_1191_),
    .A2(_1556_),
    .B1(_1557_),
    .B2(_1236_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4531_ (.A1(_1555_),
    .A2(_1558_),
    .B(_1228_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4532_ (.A1(_1416_),
    .A2(_1541_),
    .B(_1456_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4533_ (.A1(_1358_),
    .A2(_1409_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4534_ (.A1(_1407_),
    .A2(_1410_),
    .B(_1561_),
    .C(_1511_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4535_ (.A1(_1559_),
    .A2(_1560_),
    .A3(_1562_),
    .B(_1181_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4536_ (.A1(_0761_),
    .A2(_0734_),
    .A3(_0735_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4537_ (.A1(_1285_),
    .A2(_1435_),
    .A3(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4538_ (.A1(_1379_),
    .A2(_1419_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4539_ (.A1(_1130_),
    .A2(_1313_),
    .B(_1217_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4540_ (.A1(_1130_),
    .A2(_1222_),
    .B1(_1567_),
    .B2(_0735_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4541_ (.A1(_1400_),
    .A2(_1565_),
    .A3(_1566_),
    .A4(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4542_ (.A1(_1435_),
    .A2(_1564_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4543_ (.A1(_1208_),
    .A2(_1118_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4544_ (.A1(_1570_),
    .A2(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4545_ (.A1(_1563_),
    .A2(_1569_),
    .B1(_1572_),
    .B2(_1400_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4546_ (.A1(_1553_),
    .A2(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4547_ (.A1(_1323_),
    .A2(_1458_),
    .B1(_1464_),
    .B2(_1340_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4548_ (.A1(_1415_),
    .A2(_1541_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4549_ (.A1(_1273_),
    .A2(_1208_),
    .B(_1474_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4550_ (.A1(_1236_),
    .A2(_1577_),
    .B(_1454_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4551_ (.A1(_1278_),
    .A2(_1461_),
    .B1(_1544_),
    .B2(_1361_),
    .C(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4552_ (.A1(_1412_),
    .A2(_1575_),
    .B1(_1576_),
    .B2(_1456_),
    .C(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4553_ (.A1(_1433_),
    .A2(_1435_),
    .B(_1436_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4554_ (.A1(_0727_),
    .A2(_0762_),
    .A3(_0772_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4555_ (.A1(_1581_),
    .A2(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4556_ (.A1(_1278_),
    .A2(_1480_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4557_ (.A1(_1216_),
    .A2(_1142_),
    .B(_0771_),
    .C(_1180_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4558_ (.A1(_3119_),
    .A2(_1142_),
    .B(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4559_ (.A1(_1285_),
    .A2(_1583_),
    .B1(_1584_),
    .B2(_1380_),
    .C(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4560_ (.A1(_0772_),
    .A2(_1138_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4561_ (.A1(_1124_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4562_ (.A1(_1289_),
    .A2(_1583_),
    .B(_1589_),
    .C(_3131_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4563_ (.A1(_1504_),
    .A2(_1580_),
    .B(_1587_),
    .C(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4564_ (.A1(_1441_),
    .A2(_1432_),
    .A3(_1437_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4565_ (.A1(_1519_),
    .A2(_1349_),
    .A3(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4566_ (.A1(_1358_),
    .A2(_1543_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4567_ (.A1(_1373_),
    .A2(_1501_),
    .B(_1228_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4568_ (.A1(_1373_),
    .A2(_1500_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4569_ (.A1(_1110_),
    .A2(_1454_),
    .A3(_1209_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4570_ (.A1(_1453_),
    .A2(_1597_),
    .B(_1456_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4571_ (.A1(_1594_),
    .A2(_1595_),
    .B1(_1596_),
    .B2(_1185_),
    .C(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4572_ (.A1(_1518_),
    .A2(_1447_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4573_ (.A1(_1518_),
    .A2(_1447_),
    .B(_1389_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4574_ (.A1(_1339_),
    .A2(_1512_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4575_ (.I0(_1505_),
    .I1(_1602_),
    .S(_1235_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4576_ (.A1(_1440_),
    .A2(_1318_),
    .B1(_1221_),
    .B2(_0776_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4577_ (.A1(_1441_),
    .A2(_1314_),
    .B1(_1483_),
    .B2(_1603_),
    .C(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4578_ (.A1(_1469_),
    .A2(_1599_),
    .B1(_1600_),
    .B2(_1601_),
    .C(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4579_ (.A1(_1593_),
    .A2(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_1430_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4581_ (.A1(_1581_),
    .A2(_0644_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4582_ (.A1(_1608_),
    .A2(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4583_ (.A1(_1349_),
    .A2(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4584_ (.I0(_1526_),
    .I1(_1557_),
    .S(_1270_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4585_ (.I0(_0875_),
    .I1(_0951_),
    .I2(_3193_),
    .I3(_0837_),
    .S0(_1207_),
    .S1(_1269_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4586_ (.A1(_1373_),
    .A2(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4587_ (.A1(_1326_),
    .A2(_1612_),
    .B(_1614_),
    .C(_1511_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4588_ (.I(_1266_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4589_ (.A1(_1205_),
    .A2(_1616_),
    .A3(_1541_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(_1598_),
    .A2(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4591_ (.A1(_1412_),
    .A2(_1341_),
    .B(_1615_),
    .C(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4592_ (.A1(_0772_),
    .A2(_1138_),
    .B(_0770_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4593_ (.A1(_1608_),
    .A2(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4594_ (.A1(_1608_),
    .A2(_1620_),
    .B(_1389_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4595_ (.I(_1221_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4596_ (.A1(_1608_),
    .A2(_1225_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4597_ (.A1(_1140_),
    .A2(_1318_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4598_ (.A1(_1139_),
    .A2(_1623_),
    .B(_1624_),
    .C(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4599_ (.A1(_1380_),
    .A2(_1324_),
    .B1(_1621_),
    .B2(_1622_),
    .C(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4600_ (.A1(_1504_),
    .A2(_1619_),
    .B(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4601_ (.A1(_1591_),
    .A2(_1607_),
    .A3(_1611_),
    .A4(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4602_ (.A1(_1517_),
    .A2(_1537_),
    .A3(_1574_),
    .A4(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4603_ (.A1(_1427_),
    .A2(_1452_),
    .A3(_1485_),
    .A4(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4604_ (.A1(_1352_),
    .A2(_1351_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4605_ (.A1(_1351_),
    .A2(_1162_),
    .A3(_1169_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4606_ (.A1(_1387_),
    .A2(_1633_),
    .B(_1301_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4607_ (.A1(_1121_),
    .A2(_1632_),
    .B(_1634_),
    .C(_1402_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4608_ (.A1(_1405_),
    .A2(_1632_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(_1126_),
    .A2(_1315_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4610_ (.A1(_1126_),
    .A2(_1320_),
    .B(_1637_),
    .C(_1319_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_1040_),
    .A2(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4612_ (.A1(_1092_),
    .A2(_1377_),
    .A3(_1363_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4613_ (.A1(_1596_),
    .A2(_1640_),
    .B(_1367_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_1344_),
    .A2(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4615_ (.A1(_1340_),
    .A2(_1479_),
    .B1(_1505_),
    .B2(_1325_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4616_ (.A1(_1342_),
    .A2(_1509_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4617_ (.A1(_1165_),
    .A2(_1414_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4618_ (.A1(_0951_),
    .A2(_1616_),
    .B(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4619_ (.A1(_1239_),
    .A2(_1046_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4620_ (.A1(_1246_),
    .A2(_1239_),
    .B(_1647_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4621_ (.A1(_1237_),
    .A2(_1646_),
    .B1(_1648_),
    .B2(_1193_),
    .C(_1229_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4622_ (.A1(_1322_),
    .A2(_1643_),
    .B1(_1644_),
    .B2(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4623_ (.A1(_1334_),
    .A2(_1642_),
    .B1(_1650_),
    .B2(_1281_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4624_ (.A1(_1635_),
    .A2(_1636_),
    .A3(_1639_),
    .A4(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4625_ (.I(_1405_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_1147_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4627_ (.A1(_0594_),
    .A2(_1444_),
    .B(_1428_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4628_ (.A1(_1654_),
    .A2(_0505_),
    .A3(_1655_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4629_ (.A1(_0505_),
    .A2(_1655_),
    .B(_1654_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4630_ (.A1(_1656_),
    .A2(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4631_ (.A1(_1290_),
    .A2(_1656_),
    .A3(_1657_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4632_ (.A1(_1428_),
    .A2(_1449_),
    .B(_0600_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4633_ (.A1(_1654_),
    .A2(_1660_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4634_ (.A1(_1302_),
    .A2(_1661_),
    .B(_3132_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(_1342_),
    .A2(_1336_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4636_ (.A1(_1325_),
    .A2(_1613_),
    .B(_1186_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4637_ (.A1(_1198_),
    .A2(_1212_),
    .B(_1367_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4638_ (.A1(_1663_),
    .A2(_1664_),
    .B(_1665_),
    .C(_1542_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4639_ (.A1(_1158_),
    .A2(_1319_),
    .B1(_1223_),
    .B2(_1156_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4640_ (.A1(_1654_),
    .A2(_1315_),
    .B1(_1483_),
    .B2(_1279_),
    .C(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4641_ (.A1(_1469_),
    .A2(_1666_),
    .B(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4642_ (.A1(_1653_),
    .A2(_1658_),
    .B1(_1659_),
    .B2(_1662_),
    .C(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4643_ (.A1(_1392_),
    .A2(_1631_),
    .A3(_1652_),
    .A4(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4644_ (.A1(_1078_),
    .A2(_1042_),
    .A3(_1048_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4645_ (.A1(_1079_),
    .A2(_1302_),
    .A3(_1672_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4646_ (.A1(_1078_),
    .A2(_1128_),
    .A3(_1170_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4647_ (.A1(_1121_),
    .A2(_1171_),
    .A3(_1674_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4648_ (.A1(_1616_),
    .A2(_0985_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4649_ (.A1(_1080_),
    .A2(_1616_),
    .B(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4650_ (.A1(_1237_),
    .A2(_1648_),
    .B1(_1677_),
    .B2(_1193_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4651_ (.I0(_1508_),
    .I1(_1646_),
    .S(_1205_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4652_ (.A1(_1342_),
    .A2(_1679_),
    .B(_1322_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4653_ (.A1(_1367_),
    .A2(_1482_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4654_ (.A1(_1678_),
    .A2(_1680_),
    .B(_1681_),
    .C(_1331_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_1110_),
    .A2(_1202_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4656_ (.A1(_1683_),
    .A2(_1362_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4657_ (.A1(_1230_),
    .A2(_1465_),
    .B1(_1684_),
    .B2(_1301_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4658_ (.A1(_1059_),
    .A2(_1071_),
    .A3(_1073_),
    .B(_1218_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4659_ (.A1(_1076_),
    .A2(_1320_),
    .B(_1686_),
    .C(_3131_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4660_ (.A1(_1077_),
    .A2(_1225_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4661_ (.A1(_1334_),
    .A2(_1685_),
    .B(_1687_),
    .C(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4662_ (.A1(_1286_),
    .A2(_1079_),
    .A3(_1672_),
    .B(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4663_ (.A1(_3132_),
    .A2(_1673_),
    .A3(_1675_),
    .B1(_1682_),
    .B2(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4664_ (.A1(_1291_),
    .A2(_0942_),
    .A3(_0949_),
    .A4(_1295_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4665_ (.A1(_0947_),
    .A2(_1167_),
    .A3(_1304_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4666_ (.A1(_1290_),
    .A2(_1305_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4667_ (.A1(_1302_),
    .A2(_1296_),
    .A3(_1692_),
    .B1(_1693_),
    .B2(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4668_ (.A1(_1683_),
    .A2(_1415_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4669_ (.A1(_1230_),
    .A2(_1575_),
    .B1(_1696_),
    .B2(_1301_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4670_ (.A1(_1291_),
    .A2(_1315_),
    .B(_1218_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4671_ (.A1(_1291_),
    .A2(_1320_),
    .B1(_1698_),
    .B2(_1164_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4672_ (.A1(_1243_),
    .A2(_1476_),
    .B(_1412_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4673_ (.A1(_1325_),
    .A2(_1679_),
    .B(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4674_ (.A1(_1230_),
    .A2(_1584_),
    .B(_1701_),
    .C(_1331_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4675_ (.A1(_1334_),
    .A2(_1697_),
    .B(_1699_),
    .C(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4676_ (.A1(_1309_),
    .A2(_1296_),
    .A3(_1692_),
    .B(_1703_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4677_ (.A1(_1402_),
    .A2(_1695_),
    .B(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4678_ (.A1(_1691_),
    .A2(_1705_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4679_ (.A1(_1288_),
    .A2(_1348_),
    .A3(_1671_),
    .A4(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4680_ (.I(_1288_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4681_ (.A1(_3121_),
    .A2(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4682_ (.I(_1468_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4683_ (.A1(_3121_),
    .A2(_1707_),
    .B(_1709_),
    .C(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4684_ (.A1(_1708_),
    .A2(_1348_),
    .A3(_1671_),
    .A4(_1706_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4685_ (.I(_1399_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4686_ (.A1(_1713_),
    .A2(_1708_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4687_ (.A1(_3121_),
    .A2(_1712_),
    .B(_1714_),
    .C(_1317_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(_1105_),
    .A2(_1107_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4689_ (.A1(_1094_),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4690_ (.A1(_1113_),
    .A2(_1708_),
    .B(_3119_),
    .C(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4691_ (.A1(_1710_),
    .A2(_1718_),
    .A3(_1712_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4692_ (.I(_1288_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4693_ (.A1(_1113_),
    .A2(_1720_),
    .B(_1717_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4694_ (.A1(_1710_),
    .A2(_1721_),
    .B(_1312_),
    .C(_1713_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4695_ (.A1(_3119_),
    .A2(_1711_),
    .A3(_1715_),
    .B1(_1719_),
    .B2(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4696_ (.A1(_3112_),
    .A2(_3114_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4697_ (.A1(_3117_),
    .A2(_1723_),
    .B(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4698_ (.I(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4699_ (.A1(_3109_),
    .A2(_1724_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4700_ (.I(_1727_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4701_ (.A1(_1309_),
    .A2(_1553_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4702_ (.A1(_1317_),
    .A2(_1720_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4703_ (.I(_1653_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4704_ (.A1(_1317_),
    .A2(_1721_),
    .B(_1730_),
    .C(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(_1729_),
    .A2(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4706_ (.A1(\mod.pc_2[0] ),
    .A2(_0527_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4707_ (.A1(\mod.pc_2[0] ),
    .A2(_0527_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(_1727_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4709_ (.A1(_1734_),
    .A2(_1735_),
    .B(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4710_ (.A1(_1728_),
    .A2(_1733_),
    .B(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4711_ (.A1(_3105_),
    .A2(_1726_),
    .A3(_1738_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4712_ (.I(_3116_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4713_ (.A1(_1072_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4714_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4715_ (.A1(net15),
    .A2(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4716_ (.A1(net14),
    .A2(_1741_),
    .B(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4717_ (.I(\mod.ldr_hzd[12] ),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4718_ (.I(\mod.ldr_hzd[13] ),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4719_ (.I(\mod.ldr_hzd[14] ),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4720_ (.I(\mod.ldr_hzd[15] ),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4721_ (.I(_0710_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4722_ (.I(_0714_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4723_ (.I0(_1745_),
    .I1(_1746_),
    .I2(_1747_),
    .I3(_1748_),
    .S0(_1749_),
    .S1(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4724_ (.A1(_0711_),
    .A2(_0933_),
    .A3(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4725_ (.I(\mod.ldr_hzd[0] ),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4726_ (.I(\mod.ldr_hzd[1] ),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4727_ (.I(\mod.ldr_hzd[2] ),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4728_ (.I(\mod.ldr_hzd[3] ),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4729_ (.I0(_1753_),
    .I1(_1754_),
    .I2(_1755_),
    .I3(_1756_),
    .S0(_1749_),
    .S1(_1750_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4730_ (.I(\mod.ldr_hzd[9] ),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_3178_),
    .A2(_1749_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4732_ (.A1(_1758_),
    .A2(_1759_),
    .B(_3155_),
    .C(_0711_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4733_ (.I(\mod.ldr_hzd[11] ),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(_1750_),
    .A2(_3136_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4735_ (.I(\mod.ldr_hzd[10] ),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4736_ (.A1(_1761_),
    .A2(_3184_),
    .B1(_1762_),
    .B2(_1763_),
    .C1(\mod.ldr_hzd[8] ),
    .C2(_0634_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4737_ (.I(\mod.ldr_hzd[5] ),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4738_ (.A1(_1765_),
    .A2(_1759_),
    .B(_0933_),
    .C(_3147_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4739_ (.I(\mod.ldr_hzd[7] ),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4740_ (.I(\mod.ldr_hzd[6] ),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4741_ (.I(\mod.ldr_hzd[4] ),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4742_ (.A1(_1767_),
    .A2(_3184_),
    .B1(_1762_),
    .B2(_1768_),
    .C1(_1769_),
    .C2(_0634_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4743_ (.A1(_1760_),
    .A2(_1764_),
    .B1(_1766_),
    .B2(_1770_),
    .C(_0437_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4744_ (.A1(_0712_),
    .A2(_1757_),
    .B(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4745_ (.A1(_1752_),
    .A2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4746_ (.A1(_1399_),
    .A2(_1072_),
    .A3(_1740_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4747_ (.A1(_0427_),
    .A2(_0695_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4748_ (.A1(_1765_),
    .A2(_1775_),
    .B(_0693_),
    .C(_0413_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4749_ (.I(_3221_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_0613_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4751_ (.A1(_0501_),
    .A2(_0524_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4752_ (.A1(_1767_),
    .A2(_1777_),
    .B1(_1778_),
    .B2(_1769_),
    .C1(_1779_),
    .C2(_1768_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4753_ (.I(\mod.ldr_hzd[8] ),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4754_ (.A1(_1781_),
    .A2(_1778_),
    .B(_0441_),
    .C(_0657_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4755_ (.A1(\mod.ldr_hzd[11] ),
    .A2(_1777_),
    .B1(_1775_),
    .B2(\mod.ldr_hzd[9] ),
    .C1(_1779_),
    .C2(\mod.ldr_hzd[10] ),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4756_ (.A1(_1776_),
    .A2(_1780_),
    .B1(_1782_),
    .B2(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4757_ (.A1(_1748_),
    .A2(_1777_),
    .B(_0694_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4758_ (.A1(_1746_),
    .A2(_1775_),
    .B1(_1778_),
    .B2(_1745_),
    .C1(_1779_),
    .C2(_1747_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4759_ (.A1(_1785_),
    .A2(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4760_ (.A1(_0657_),
    .A2(_0693_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1754_),
    .A2(_1775_),
    .B(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4762_ (.A1(_1756_),
    .A2(_1777_),
    .B1(_1778_),
    .B2(_1753_),
    .C1(_1779_),
    .C2(_1755_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4763_ (.A1(_1789_),
    .A2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4764_ (.A1(_1784_),
    .A2(_1787_),
    .A3(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(\mod.instr_2[4] ),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4766_ (.I(_0523_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4767_ (.A1(_1793_),
    .A2(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4768_ (.I(_1795_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4769_ (.I(_1793_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4770_ (.A1(_1797_),
    .A2(_1794_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4772_ (.A1(\mod.ldr_hzd[1] ),
    .A2(_1796_),
    .B1(_1799_),
    .B2(\mod.ldr_hzd[3] ),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4773_ (.A1(_1797_),
    .A2(\mod.instr_2[3] ),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4774_ (.I(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_1793_),
    .A2(\mod.instr_2[3] ),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4776_ (.I(\mod.instr_2[5] ),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4777_ (.A1(\mod.ldr_hzd[2] ),
    .A2(_1802_),
    .B1(_1803_),
    .B2(\mod.ldr_hzd[0] ),
    .C(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(\mod.ldr_hzd[5] ),
    .A2(_1796_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4779_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_1801_),
    .B1(_1803_),
    .B2(\mod.ldr_hzd[4] ),
    .C1(_1798_),
    .C2(\mod.ldr_hzd[7] ),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4780_ (.A1(\mod.instr_2[5] ),
    .A2(_1806_),
    .A3(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(\mod.instr_2[6] ),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4782_ (.A1(_1800_),
    .A2(_1805_),
    .B(_1808_),
    .C(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4783_ (.A1(_1758_),
    .A2(_1796_),
    .B1(_1799_),
    .B2(_1761_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4784_ (.I(_1803_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4785_ (.A1(_1763_),
    .A2(_1802_),
    .B1(_1812_),
    .B2(_1781_),
    .C(_1804_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4786_ (.A1(\mod.ldr_hzd[14] ),
    .A2(_1802_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4787_ (.A1(\mod.ldr_hzd[13] ),
    .A2(_1795_),
    .B1(_1803_),
    .B2(\mod.ldr_hzd[12] ),
    .C1(_1799_),
    .C2(\mod.ldr_hzd[15] ),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4788_ (.A1(_1804_),
    .A2(_1814_),
    .A3(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4789_ (.A1(\mod.instr_2[6] ),
    .A2(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4790_ (.A1(_1811_),
    .A2(_1813_),
    .B(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4791_ (.A1(_1810_),
    .A2(_1818_),
    .B(_1774_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4792_ (.A1(_1774_),
    .A2(_1792_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4793_ (.A1(_1767_),
    .A2(_1768_),
    .A3(_1765_),
    .A4(_1769_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4794_ (.A1(_1761_),
    .A2(_1763_),
    .A3(_1758_),
    .A4(_1781_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4795_ (.A1(_1748_),
    .A2(_1747_),
    .A3(_1746_),
    .A4(_1745_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4796_ (.A1(_1756_),
    .A2(_1755_),
    .A3(_1754_),
    .A4(_1753_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4797_ (.A1(_1822_),
    .A2(_1823_),
    .A3(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4798_ (.A1(_1773_),
    .A2(_1820_),
    .B1(_1821_),
    .B2(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4799_ (.A1(_1744_),
    .A2(_1826_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4800_ (.I(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(_1725_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4802_ (.A1(\mod.valid2 ),
    .A2(_1827_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4803_ (.I(net13),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4804_ (.A1(_1829_),
    .A2(_1830_),
    .B(\mod.valid0 ),
    .C(_1831_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4805_ (.A1(_1828_),
    .A2(_1832_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4806_ (.I(_1833_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4807_ (.I(_1834_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_3104_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4809_ (.I(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4810_ (.I(_1725_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4811_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4812_ (.A1(_1837_),
    .A2(_1839_),
    .B(\mod.pc[0] ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4813_ (.I(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4814_ (.A1(_1836_),
    .A2(_1838_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4815_ (.I(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4816_ (.A1(_1843_),
    .A2(_1833_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4817_ (.I(_1844_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4818_ (.A1(\mod.pc0[0] ),
    .A2(_1835_),
    .B1(_1841_),
    .B2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4819_ (.A1(_1739_),
    .A2(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4820_ (.I(_3097_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4821_ (.I(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4822_ (.A1(_0738_),
    .A2(_0746_),
    .B(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4823_ (.I(_3093_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4824_ (.I(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(_1848_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4826_ (.A1(_1853_),
    .A2(_1733_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4827_ (.A1(_3102_),
    .A2(_1847_),
    .B1(_1850_),
    .B2(_1852_),
    .C(_1854_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(_1836_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4829_ (.A1(_1855_),
    .A2(_1829_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4831_ (.I(_1309_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(_1858_),
    .A2(_1573_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_1072_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(_3111_),
    .A2(_3115_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4835_ (.A1(_1860_),
    .A2(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4836_ (.A1(_0730_),
    .A2(_0503_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4837_ (.A1(_1735_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4838_ (.A1(_1862_),
    .A2(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4839_ (.A1(_1728_),
    .A2(_1859_),
    .B(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4840_ (.I(\mod.pc0[1] ),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4841_ (.I(_1843_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4842_ (.A1(\mod.pc[1] ),
    .A2(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4843_ (.A1(_1867_),
    .A2(_1835_),
    .B1(_1845_),
    .B2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4844_ (.A1(_1857_),
    .A2(_1866_),
    .B(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4845_ (.A1(_0689_),
    .A2(_0702_),
    .B(_1849_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4846_ (.I(_1858_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4847_ (.A1(_1873_),
    .A2(_1573_),
    .B(_3098_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4848_ (.A1(_3102_),
    .A2(_1871_),
    .B1(_1872_),
    .B2(_1852_),
    .C(_1874_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(\mod.des.des_counter[0] ),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4850_ (.I(_1875_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4851_ (.A1(_1653_),
    .A2(_1591_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4852_ (.A1(_0608_),
    .A2(_0618_),
    .B(_1849_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4853_ (.I(_1862_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4854_ (.I(_0447_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4855_ (.A1(_0730_),
    .A2(_0503_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4856_ (.A1(_1735_),
    .A2(_1863_),
    .B(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4857_ (.A1(_0622_),
    .A2(_1880_),
    .A3(_1882_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_1862_),
    .A2(_1877_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4859_ (.A1(_1879_),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4860_ (.A1(_3105_),
    .A2(_1838_),
    .A3(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(_1834_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4862_ (.I(\mod.pc[2] ),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4863_ (.I(_1833_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4864_ (.I(_1842_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4865_ (.I(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4867_ (.A1(_1888_),
    .A2(_1889_),
    .B(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4868_ (.A1(\mod.pc0[2] ),
    .A2(_1887_),
    .B(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4869_ (.A1(_3101_),
    .A2(_1886_),
    .A3(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4870_ (.A1(_1876_),
    .A2(_1877_),
    .B1(_1878_),
    .B2(_1852_),
    .C(_1895_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4871_ (.A1(_1611_),
    .A2(_1628_),
    .B(_1731_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4872_ (.I(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4873_ (.A1(_0000_),
    .A2(_0675_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4874_ (.I(_3099_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4875_ (.I(_1727_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4876_ (.I(_0830_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4877_ (.A1(_0766_),
    .A2(_1880_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4878_ (.A1(_0766_),
    .A2(_1880_),
    .B1(_1735_),
    .B2(_1863_),
    .C(_1881_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4879_ (.A1(_1902_),
    .A2(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4880_ (.A1(_0676_),
    .A2(_1901_),
    .A3(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_1736_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4882_ (.A1(_1900_),
    .A2(_1896_),
    .B(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4883_ (.A1(_3105_),
    .A2(_1726_),
    .A3(_1907_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_1834_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4885_ (.A1(_1837_),
    .A2(_1839_),
    .B(\mod.pc[3] ),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4886_ (.I(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4887_ (.A1(\mod.pc0[3] ),
    .A2(_1909_),
    .B1(_1845_),
    .B2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4888_ (.A1(_1899_),
    .A2(_1908_),
    .A3(_1912_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4889_ (.A1(_1876_),
    .A2(_1897_),
    .B1(_1898_),
    .B2(_1852_),
    .C(_1913_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4890_ (.A1(_1653_),
    .A2(_1607_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(_1848_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4892_ (.A1(_0553_),
    .A2(_0561_),
    .B(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4893_ (.I(_3094_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4894_ (.I(\mod.pc_2[4] ),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_0871_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4896_ (.A1(\mod.pc_2[3] ),
    .A2(_1901_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(\mod.pc_2[3] ),
    .A2(_1901_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4898_ (.A1(_1902_),
    .A2(_1920_),
    .A3(_1903_),
    .B(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4899_ (.A1(_1918_),
    .A2(_1919_),
    .A3(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4900_ (.A1(_1736_),
    .A2(_1914_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4901_ (.A1(_1728_),
    .A2(_1923_),
    .B(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4902_ (.A1(_3105_),
    .A2(_1726_),
    .A3(_1925_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4903_ (.I(\mod.pc[4] ),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(_1833_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4905_ (.A1(_1927_),
    .A2(_1928_),
    .B(_1892_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4906_ (.A1(\mod.pc0[4] ),
    .A2(_1887_),
    .B(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4907_ (.A1(_1899_),
    .A2(_1926_),
    .A3(_1930_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4908_ (.A1(_1876_),
    .A2(_1914_),
    .B1(_1916_),
    .B2(_1917_),
    .C(_1931_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4909_ (.I(_1736_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4910_ (.A1(_1858_),
    .A2(_1537_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4911_ (.I(_0935_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4912_ (.A1(_1918_),
    .A2(_1919_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4913_ (.A1(_1918_),
    .A2(_1919_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4914_ (.A1(_1935_),
    .A2(_1922_),
    .B(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4915_ (.A1(_0506_),
    .A2(_1934_),
    .A3(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4916_ (.A1(_1900_),
    .A2(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4917_ (.A1(_1932_),
    .A2(_1933_),
    .B(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4918_ (.A1(_1855_),
    .A2(_1726_),
    .A3(_1940_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4919_ (.I(_1836_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4920_ (.I(_1838_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4921_ (.A1(_1942_),
    .A2(_1943_),
    .B(\mod.pc[5] ),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4922_ (.I(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4923_ (.A1(\mod.pc0[5] ),
    .A2(_1835_),
    .B1(_1845_),
    .B2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4924_ (.A1(_1941_),
    .A2(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4925_ (.A1(_0532_),
    .A2(_0536_),
    .B(_3092_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4926_ (.I(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4927_ (.A1(_3098_),
    .A2(_1933_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4928_ (.A1(_3102_),
    .A2(_1947_),
    .B1(_1949_),
    .B2(_1917_),
    .C(_1950_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4929_ (.A1(_1452_),
    .A2(_1485_),
    .B(_1858_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4930_ (.A1(_0486_),
    .A2(_0496_),
    .B(_1915_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(_0903_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(_0506_),
    .A2(_1934_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4933_ (.A1(_1954_),
    .A2(_1937_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4934_ (.A1(_0506_),
    .A2(_1934_),
    .B(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4935_ (.A1(_0453_),
    .A2(_1953_),
    .A3(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4936_ (.A1(_1862_),
    .A2(_1951_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4937_ (.A1(_1879_),
    .A2(_1957_),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4938_ (.A1(_1837_),
    .A2(_1839_),
    .A3(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_1844_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4940_ (.A1(_1942_),
    .A2(_1943_),
    .B(\mod.pc[6] ),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4941_ (.I(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4942_ (.A1(\mod.pc0[6] ),
    .A2(_1909_),
    .B1(_1961_),
    .B2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4943_ (.A1(_1899_),
    .A2(_1960_),
    .A3(_1964_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4944_ (.A1(_1876_),
    .A2(_1951_),
    .B1(_1952_),
    .B2(_1917_),
    .C(_1965_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4945_ (.I(_1875_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4946_ (.A1(_1731_),
    .A2(_1670_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4947_ (.I(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4948_ (.A1(_0411_),
    .A2(_0433_),
    .B(_1915_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4949_ (.I(_1036_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4950_ (.A1(_0452_),
    .A2(_1953_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4951_ (.A1(_0452_),
    .A2(_1953_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4952_ (.A1(_1971_),
    .A2(_1956_),
    .B(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4953_ (.A1(_0596_),
    .A2(_1970_),
    .A3(_1973_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4954_ (.A1(_1900_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4955_ (.A1(_1932_),
    .A2(_1967_),
    .B(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4956_ (.A1(_1855_),
    .A2(_1829_),
    .A3(_1976_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4957_ (.A1(_1942_),
    .A2(_1943_),
    .B(\mod.pc[7] ),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4958_ (.I(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4959_ (.A1(\mod.pc0[7] ),
    .A2(_1909_),
    .B1(_1961_),
    .B2(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4960_ (.A1(_1899_),
    .A2(_1977_),
    .A3(_1980_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4961_ (.A1(_1966_),
    .A2(_1968_),
    .B1(_1969_),
    .B2(_1917_),
    .C(_1981_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4962_ (.I(\mod.pc[8] ),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4963_ (.A1(_1982_),
    .A2(_1889_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4964_ (.A1(\mod.pc0[8] ),
    .A2(_1835_),
    .B(_1983_),
    .C(_1857_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4965_ (.I(_1728_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4966_ (.A1(_1873_),
    .A2(_1517_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4967_ (.I(_1004_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4968_ (.A1(\mod.pc_2[7] ),
    .A2(_1970_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4969_ (.A1(\mod.pc_2[7] ),
    .A2(_1970_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4970_ (.A1(_1988_),
    .A2(_1973_),
    .B(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4971_ (.A1(_0779_),
    .A2(_1987_),
    .A3(_1990_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4972_ (.A1(_1932_),
    .A2(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4973_ (.A1(_1985_),
    .A2(_1986_),
    .B(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4974_ (.A1(_1891_),
    .A2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4975_ (.A1(_1984_),
    .A2(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4976_ (.A1(_0815_),
    .A2(_0826_),
    .B(_1915_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4977_ (.I(_3094_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4978_ (.A1(_1873_),
    .A2(_1517_),
    .B(_3098_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4979_ (.A1(_3101_),
    .A2(_1995_),
    .B1(_1996_),
    .B2(_1997_),
    .C(_1998_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4980_ (.A1(_1873_),
    .A2(_1427_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4981_ (.A1(_0861_),
    .A2(_0867_),
    .B(_1853_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4982_ (.I(_1843_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4983_ (.A1(_0833_),
    .A2(_1987_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(_0833_),
    .A2(_1987_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4985_ (.A1(_2002_),
    .A2(_1990_),
    .B(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4986_ (.I(\mod.pc_2[9] ),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4987_ (.A1(_0441_),
    .A2(_1034_),
    .B(_1035_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4988_ (.A1(_2005_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4989_ (.A1(_2005_),
    .A2(_2006_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4990_ (.A1(_2007_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4991_ (.A1(_2004_),
    .A2(_2009_),
    .B(_1900_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4992_ (.A1(_2004_),
    .A2(_2009_),
    .B(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4993_ (.A1(_1879_),
    .A2(_1999_),
    .B(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4994_ (.A1(_2001_),
    .A2(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4995_ (.I(\mod.pc[9] ),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4996_ (.A1(_2014_),
    .A2(_1928_),
    .B(_1892_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4997_ (.A1(\mod.pc0[9] ),
    .A2(_1887_),
    .B(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4998_ (.A1(_3100_),
    .A2(_2013_),
    .A3(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4999_ (.A1(_1966_),
    .A2(_1999_),
    .B1(_2000_),
    .B2(_1997_),
    .C(_2017_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5000_ (.A1(\mod.pc0[10] ),
    .A2(_1889_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5001_ (.I(\mod.pc[10] ),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5002_ (.A1(_2019_),
    .A2(_1887_),
    .B(_2001_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5003_ (.I(_1731_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5004_ (.A1(_2021_),
    .A2(_1705_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5005_ (.A1(_2004_),
    .A2(_2008_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5006_ (.A1(_0911_),
    .A2(_1106_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5007_ (.A1(_2007_),
    .A2(_2023_),
    .A3(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(_2024_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5009_ (.A1(_2007_),
    .A2(_2023_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5010_ (.A1(_2026_),
    .A2(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5011_ (.A1(_1932_),
    .A2(_2025_),
    .A3(_2028_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5012_ (.A1(_1985_),
    .A2(_2022_),
    .B(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5013_ (.A1(_2018_),
    .A2(_2020_),
    .B1(_2030_),
    .B2(_2001_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5014_ (.A1(_0926_),
    .A2(_0930_),
    .B(_1853_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5015_ (.A1(_3092_),
    .A2(_2022_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5016_ (.A1(_3101_),
    .A2(_2031_),
    .B1(_2032_),
    .B2(_1997_),
    .C(_2033_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5017_ (.A1(_2021_),
    .A2(_1348_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5018_ (.A1(_0895_),
    .A2(_0900_),
    .B(_1853_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5019_ (.I0(\mod.pc0[11] ),
    .I1(\mod.pc[11] ),
    .S(_1834_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5020_ (.I(_1879_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5021_ (.A1(\mod.pc_2[10] ),
    .A2(_1106_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5022_ (.A1(_2038_),
    .A2(_2028_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5023_ (.A1(_0563_),
    .A2(_1034_),
    .B(_1035_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5024_ (.A1(_0878_),
    .A2(_2040_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5025_ (.A1(_2039_),
    .A2(_2041_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5026_ (.A1(_2037_),
    .A2(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5027_ (.A1(_2037_),
    .A2(_2034_),
    .B(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5028_ (.I0(_2036_),
    .I1(_2044_),
    .S(_2001_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5029_ (.A1(_1875_),
    .A2(_3094_),
    .A3(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5030_ (.A1(_1966_),
    .A2(_2034_),
    .B1(_2035_),
    .B2(_1997_),
    .C(_2046_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5031_ (.A1(_2021_),
    .A2(_1652_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5032_ (.I(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5033_ (.A1(_0000_),
    .A2(_1032_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5034_ (.A1(\mod.pc_2[11] ),
    .A2(_2040_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5035_ (.A1(_2039_),
    .A2(_2041_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5036_ (.A1(\mod.pc_2[12] ),
    .A2(_1074_),
    .A3(_2051_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_1985_),
    .A2(_2052_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5038_ (.A1(_1985_),
    .A2(_2047_),
    .B(_2053_),
    .C(_1843_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5039_ (.I(\mod.pc[12] ),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5040_ (.A1(_2055_),
    .A2(_1928_),
    .B(_1892_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5041_ (.A1(\mod.pc0[12] ),
    .A2(_1909_),
    .B(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5042_ (.A1(_3100_),
    .A2(_2054_),
    .A3(_2057_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5043_ (.A1(_1966_),
    .A2(_2048_),
    .B1(_2049_),
    .B2(_1851_),
    .C(_2058_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(_2021_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5045_ (.A1(_2059_),
    .A2(_1392_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5046_ (.A1(_1849_),
    .A2(_1001_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5047_ (.I(_1044_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_2062_),
    .A2(_1074_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5049_ (.A1(_2062_),
    .A2(_1074_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5050_ (.A1(_2063_),
    .A2(_2051_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5051_ (.A1(_0957_),
    .A2(\mod.funct7[2] ),
    .A3(_2065_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5052_ (.A1(_2037_),
    .A2(_2060_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5053_ (.A1(_2037_),
    .A2(_2066_),
    .B(_2067_),
    .C(_1868_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5054_ (.I(\mod.pc[13] ),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5055_ (.A1(_2069_),
    .A2(_1868_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5056_ (.A1(\mod.pc0[13] ),
    .A2(_1889_),
    .B1(_1961_),
    .B2(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5057_ (.A1(_3100_),
    .A2(_2068_),
    .A3(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5058_ (.A1(_1875_),
    .A2(_2060_),
    .B1(_2061_),
    .B2(_1851_),
    .C(_2072_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5059_ (.A1(_2059_),
    .A2(_1691_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5060_ (.A1(_3097_),
    .A2(_3093_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5061_ (.A1(_0000_),
    .A2(_1851_),
    .A3(_1069_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5062_ (.A1(_2073_),
    .A2(_2074_),
    .B(_2075_),
    .ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5063_ (.A1(_1848_),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5064_ (.A1(_2059_),
    .A2(_1720_),
    .A3(_2074_),
    .B1(_2076_),
    .B2(_1103_),
    .ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5065_ (.A1(_1860_),
    .A2(_1740_),
    .A3(_1830_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5066_ (.I(_2077_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5067_ (.A1(_1713_),
    .A2(net22),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5068_ (.I(_2078_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5069_ (.I(net11),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_2079_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5071_ (.I(_2080_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5072_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5074_ (.I(_2081_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5075_ (.A1(\mod.rd_3[2] ),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5076_ (.A1(_0440_),
    .A2(_2082_),
    .B(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5077_ (.I(_1809_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5078_ (.I(_2081_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5079_ (.A1(\mod.rd_3[3] ),
    .A2(_2083_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5080_ (.A1(_2086_),
    .A2(_2087_),
    .B(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5081_ (.A1(_2085_),
    .A2(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(net12),
    .A2(_2082_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5083_ (.I(\mod.valid2 ),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5084_ (.A1(net12),
    .A2(_1828_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5085_ (.A1(_2092_),
    .A2(_1740_),
    .A3(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5086_ (.A1(\mod.rd_3[1] ),
    .A2(_2083_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5087_ (.A1(_1797_),
    .A2(_2082_),
    .B(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5088_ (.A1(_2091_),
    .A2(_2094_),
    .B(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5089_ (.A1(\mod.rd_3[0] ),
    .A2(_2083_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5090_ (.A1(_1794_),
    .A2(_2082_),
    .B(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5091_ (.A1(_2097_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5092_ (.A1(_2090_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5093_ (.I(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(_2102_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_2087_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_1724_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(_2106_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5099_ (.I(_2106_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5100_ (.A1(_2108_),
    .A2(_1733_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5101_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(_1860_),
    .A2(_3124_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5103_ (.A1(_2110_),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5104_ (.I(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5105_ (.A1(_1133_),
    .A2(_2107_),
    .B(_2109_),
    .C(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5106_ (.A1(\mod.des.des_dout[21] ),
    .A2(_2105_),
    .B(_2114_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5107_ (.I(_2115_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5108_ (.I(_2101_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5109_ (.I(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5110_ (.A1(\mod.registers.r1[0] ),
    .A2(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5111_ (.A1(_2103_),
    .A2(_2116_),
    .B(_2119_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_1861_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5113_ (.I(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5114_ (.I(_2112_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5115_ (.I(_1861_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5116_ (.A1(_0730_),
    .A2(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5117_ (.A1(_2121_),
    .A2(_1859_),
    .B(_2122_),
    .C(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5118_ (.A1(\mod.des.des_dout[22] ),
    .A2(_2105_),
    .B(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5119_ (.I(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5120_ (.A1(\mod.registers.r1[1] ),
    .A2(_2118_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5121_ (.A1(_2103_),
    .A2(_2127_),
    .B(_2128_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5122_ (.I(_2120_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5123_ (.A1(_0766_),
    .A2(_2123_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5124_ (.A1(_2129_),
    .A2(_1877_),
    .B(_2122_),
    .C(_2130_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5125_ (.A1(\mod.des.des_dout[23] ),
    .A2(_2105_),
    .B(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5126_ (.I(_2132_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5127_ (.A1(\mod.registers.r1[2] ),
    .A2(_2118_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5128_ (.A1(_2103_),
    .A2(_2133_),
    .B(_2134_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5129_ (.A1(_2108_),
    .A2(_1896_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5130_ (.A1(_0676_),
    .A2(_2107_),
    .B(_2122_),
    .C(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5131_ (.A1(\mod.des.des_dout[24] ),
    .A2(_2105_),
    .B(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5132_ (.I(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5133_ (.A1(\mod.registers.r1[3] ),
    .A2(_2118_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5134_ (.A1(_2103_),
    .A2(_2138_),
    .B(_2139_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5135_ (.I(_2102_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5136_ (.I(_2104_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5137_ (.A1(_1918_),
    .A2(_2120_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5138_ (.A1(_2129_),
    .A2(_1914_),
    .B(_2122_),
    .C(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5139_ (.A1(\mod.des.des_dout[25] ),
    .A2(_2141_),
    .B(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5140_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5141_ (.I(_2117_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5142_ (.A1(\mod.registers.r1[4] ),
    .A2(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5143_ (.A1(_2140_),
    .A2(_2145_),
    .B(_2147_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5144_ (.I(_2111_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5145_ (.I(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5146_ (.A1(_2129_),
    .A2(_1933_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5147_ (.A1(_0591_),
    .A2(_2121_),
    .B(_2149_),
    .C(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5148_ (.I(_2087_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5149_ (.I(_2111_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5150_ (.A1(_0527_),
    .A2(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5151_ (.A1(_2152_),
    .A2(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5152_ (.A1(\mod.des.des_dout[26] ),
    .A2(_2141_),
    .B1(_2151_),
    .B2(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5153_ (.I(_2156_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5154_ (.A1(\mod.registers.r1[5] ),
    .A2(_2146_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5155_ (.A1(_2140_),
    .A2(_2157_),
    .B(_2158_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5156_ (.I(_2110_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(_2120_),
    .A2(_1951_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5158_ (.A1(_0452_),
    .A2(_2129_),
    .B(_2148_),
    .C(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5159_ (.A1(_3109_),
    .A2(_3165_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5160_ (.I(_2162_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(_0503_),
    .A2(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5162_ (.A1(_2159_),
    .A2(_2161_),
    .A3(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5163_ (.A1(\mod.des.des_dout[27] ),
    .A2(_2159_),
    .B(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5164_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5165_ (.A1(\mod.registers.r1[6] ),
    .A2(_2146_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5166_ (.A1(_2140_),
    .A2(_2167_),
    .B(_2168_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5167_ (.A1(_2123_),
    .A2(_1967_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5168_ (.A1(_0596_),
    .A2(_2121_),
    .B(_2149_),
    .C(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5169_ (.A1(_1880_),
    .A2(_2153_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5170_ (.A1(_2152_),
    .A2(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5171_ (.A1(\mod.des.des_dout[28] ),
    .A2(_2141_),
    .B1(_2170_),
    .B2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5172_ (.I(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5173_ (.A1(\mod.registers.r1[7] ),
    .A2(_2146_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5174_ (.A1(_2140_),
    .A2(_2174_),
    .B(_2175_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5175_ (.I(_2102_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5176_ (.I(_2106_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5177_ (.I(_2106_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5178_ (.A1(_0833_),
    .A2(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5179_ (.A1(_2177_),
    .A2(_1986_),
    .B(_2149_),
    .C(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5180_ (.A1(_1901_),
    .A2(_2153_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5181_ (.A1(_2152_),
    .A2(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5182_ (.A1(\mod.des.des_dout[29] ),
    .A2(_2141_),
    .B1(_2180_),
    .B2(_2182_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5183_ (.I(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5184_ (.I(_2117_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5185_ (.A1(\mod.registers.r1[8] ),
    .A2(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5186_ (.A1(_2176_),
    .A2(_2184_),
    .B(_2186_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5187_ (.I(_2087_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_2005_),
    .A2(_2178_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5189_ (.A1(_2177_),
    .A2(_1999_),
    .B(_2149_),
    .C(_2188_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5190_ (.I(_2110_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(_1919_),
    .A2(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_2113_),
    .A2(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5193_ (.A1(\mod.des.des_dout[30] ),
    .A2(_2187_),
    .B1(_2189_),
    .B2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5194_ (.I(_2193_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5195_ (.A1(\mod.registers.r1[9] ),
    .A2(_2185_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5196_ (.A1(_2176_),
    .A2(_2194_),
    .B(_2195_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5197_ (.I(_2148_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5198_ (.A1(\mod.pc_2[10] ),
    .A2(_2178_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5199_ (.A1(_2177_),
    .A2(_2022_),
    .B(_2196_),
    .C(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5200_ (.A1(_1934_),
    .A2(_2153_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5201_ (.A1(_2104_),
    .A2(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5202_ (.A1(\mod.des.des_dout[31] ),
    .A2(_2187_),
    .B1(_2198_),
    .B2(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5203_ (.I(_2201_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5204_ (.A1(\mod.registers.r1[10] ),
    .A2(_2185_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5205_ (.A1(_2176_),
    .A2(_2202_),
    .B(_2203_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(\mod.pc_2[11] ),
    .A2(_2108_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5207_ (.A1(_2177_),
    .A2(_2034_),
    .B(_2196_),
    .C(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5208_ (.A1(_1953_),
    .A2(_2148_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5209_ (.A1(_2104_),
    .A2(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5210_ (.A1(\mod.des.des_dout[32] ),
    .A2(_2187_),
    .B1(_2205_),
    .B2(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5211_ (.I(_2208_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5212_ (.A1(\mod.registers.r1[11] ),
    .A2(_2185_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5213_ (.A1(_2176_),
    .A2(_2209_),
    .B(_2210_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5214_ (.I(_2102_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5215_ (.A1(_2123_),
    .A2(_2047_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5216_ (.A1(_2062_),
    .A2(_2121_),
    .B(_2196_),
    .C(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5217_ (.A1(_1970_),
    .A2(_2190_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5218_ (.A1(_2113_),
    .A2(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5219_ (.A1(\mod.des.des_dout[33] ),
    .A2(_2187_),
    .B1(_2213_),
    .B2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5220_ (.I(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5221_ (.I(_2117_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(\mod.registers.r1[12] ),
    .A2(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5223_ (.A1(_2211_),
    .A2(_2217_),
    .B(_2219_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5224_ (.A1(\mod.pc_2[13] ),
    .A2(_2108_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5225_ (.A1(_2107_),
    .A2(_2060_),
    .B(_2196_),
    .C(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5226_ (.A1(_1987_),
    .A2(_2110_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5227_ (.A1(_2113_),
    .A2(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5228_ (.A1(\mod.des.des_dout[34] ),
    .A2(_2152_),
    .B1(_2221_),
    .B2(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5229_ (.I(_2224_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5230_ (.A1(\mod.registers.r1[13] ),
    .A2(_2218_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5231_ (.A1(_2211_),
    .A2(_2225_),
    .B(_2226_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5232_ (.A1(_2107_),
    .A2(_2073_),
    .A3(_2163_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5233_ (.A1(_2006_),
    .A2(_2163_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(_2190_),
    .A2(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5235_ (.A1(\mod.des.des_dout[35] ),
    .A2(_2159_),
    .B1(_2227_),
    .B2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5236_ (.I(_2230_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(\mod.registers.r1[14] ),
    .A2(_2218_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(_2211_),
    .A2(_2231_),
    .B(_2232_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5239_ (.A1(_2178_),
    .A2(_2059_),
    .A3(_1720_),
    .A4(_2163_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5240_ (.A1(_1106_),
    .A2(_2162_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5241_ (.A1(_2190_),
    .A2(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5242_ (.A1(\mod.des.des_dout[36] ),
    .A2(_2159_),
    .B1(_2233_),
    .B2(_2235_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5243_ (.I(_2236_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(\mod.registers.r1[15] ),
    .A2(_2218_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5245_ (.A1(_2211_),
    .A2(_2237_),
    .B(_2238_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5246_ (.A1(_2091_),
    .A2(_2094_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5247_ (.A1(_2239_),
    .A2(_2096_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5248_ (.A1(_2099_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(_2090_),
    .A2(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5250_ (.I(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5252_ (.I(_2242_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5253_ (.I(_2245_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(\mod.registers.r2[0] ),
    .A2(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5255_ (.A1(_2116_),
    .A2(_2244_),
    .B(_2247_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5256_ (.A1(\mod.registers.r2[1] ),
    .A2(_2246_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5257_ (.A1(_2127_),
    .A2(_2244_),
    .B(_2248_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(\mod.registers.r2[2] ),
    .A2(_2246_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5259_ (.A1(_2133_),
    .A2(_2244_),
    .B(_2249_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5260_ (.A1(\mod.registers.r2[3] ),
    .A2(_2246_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5261_ (.A1(_2138_),
    .A2(_2244_),
    .B(_2250_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5262_ (.I(_2243_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5263_ (.I(_2245_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5264_ (.A1(\mod.registers.r2[4] ),
    .A2(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5265_ (.A1(_2145_),
    .A2(_2251_),
    .B(_2253_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(\mod.registers.r2[5] ),
    .A2(_2252_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5267_ (.A1(_2157_),
    .A2(_2251_),
    .B(_2254_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(\mod.registers.r2[6] ),
    .A2(_2252_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5269_ (.A1(_2167_),
    .A2(_2251_),
    .B(_2255_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5270_ (.A1(\mod.registers.r2[7] ),
    .A2(_2252_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5271_ (.A1(_2174_),
    .A2(_2251_),
    .B(_2256_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5272_ (.I(_2243_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5273_ (.I(_2245_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(\mod.registers.r2[8] ),
    .A2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5275_ (.A1(_2184_),
    .A2(_2257_),
    .B(_2259_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5276_ (.A1(\mod.registers.r2[9] ),
    .A2(_2258_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5277_ (.A1(_2194_),
    .A2(_2257_),
    .B(_2260_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(\mod.registers.r2[10] ),
    .A2(_2258_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5279_ (.A1(_2202_),
    .A2(_2257_),
    .B(_2261_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5280_ (.A1(\mod.registers.r2[11] ),
    .A2(_2258_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5281_ (.A1(_2209_),
    .A2(_2257_),
    .B(_2262_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5282_ (.I(_2243_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5283_ (.I(_2245_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(\mod.registers.r2[12] ),
    .A2(_2264_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5285_ (.A1(_2217_),
    .A2(_2263_),
    .B(_2265_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5286_ (.A1(\mod.registers.r2[13] ),
    .A2(_2264_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5287_ (.A1(_2225_),
    .A2(_2263_),
    .B(_2266_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5288_ (.A1(\mod.registers.r2[14] ),
    .A2(_2264_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5289_ (.A1(_2231_),
    .A2(_2263_),
    .B(_2267_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5290_ (.A1(\mod.registers.r2[15] ),
    .A2(_2264_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5291_ (.A1(_2237_),
    .A2(_2263_),
    .B(_2268_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5292_ (.I(_2099_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5293_ (.A1(_2269_),
    .A2(_2240_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5294_ (.A1(_2090_),
    .A2(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5295_ (.I(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5296_ (.I(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5297_ (.I(_2271_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5298_ (.I(_2274_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(\mod.registers.r3[0] ),
    .A2(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5300_ (.A1(_2116_),
    .A2(_2273_),
    .B(_2276_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5301_ (.A1(\mod.registers.r3[1] ),
    .A2(_2275_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5302_ (.A1(_2127_),
    .A2(_2273_),
    .B(_2277_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5303_ (.A1(\mod.registers.r3[2] ),
    .A2(_2275_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5304_ (.A1(_2133_),
    .A2(_2273_),
    .B(_2278_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5305_ (.A1(\mod.registers.r3[3] ),
    .A2(_2275_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5306_ (.A1(_2138_),
    .A2(_2273_),
    .B(_2279_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5307_ (.I(_2272_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5308_ (.I(_2274_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5309_ (.A1(\mod.registers.r3[4] ),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5310_ (.A1(_2145_),
    .A2(_2280_),
    .B(_2282_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5311_ (.A1(\mod.registers.r3[5] ),
    .A2(_2281_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5312_ (.A1(_2157_),
    .A2(_2280_),
    .B(_2283_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5313_ (.A1(\mod.registers.r3[6] ),
    .A2(_2281_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5314_ (.A1(_2167_),
    .A2(_2280_),
    .B(_2284_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5315_ (.A1(\mod.registers.r3[7] ),
    .A2(_2281_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5316_ (.A1(_2174_),
    .A2(_2280_),
    .B(_2285_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5317_ (.I(_2272_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5318_ (.I(_2274_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(\mod.registers.r3[8] ),
    .A2(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5320_ (.A1(_2184_),
    .A2(_2286_),
    .B(_2288_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5321_ (.A1(\mod.registers.r3[9] ),
    .A2(_2287_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5322_ (.A1(_2194_),
    .A2(_2286_),
    .B(_2289_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5323_ (.A1(\mod.registers.r3[10] ),
    .A2(_2287_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5324_ (.A1(_2202_),
    .A2(_2286_),
    .B(_2290_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5325_ (.A1(\mod.registers.r3[11] ),
    .A2(_2287_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5326_ (.A1(_2209_),
    .A2(_2286_),
    .B(_2291_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5327_ (.I(_2272_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_2274_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5329_ (.A1(\mod.registers.r3[12] ),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5330_ (.A1(_2217_),
    .A2(_2292_),
    .B(_2294_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5331_ (.A1(\mod.registers.r3[13] ),
    .A2(_2293_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5332_ (.A1(_2225_),
    .A2(_2292_),
    .B(_2295_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(\mod.registers.r3[14] ),
    .A2(_2293_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5334_ (.A1(_2231_),
    .A2(_2292_),
    .B(_2296_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5335_ (.A1(\mod.registers.r3[15] ),
    .A2(_2293_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5336_ (.A1(_2237_),
    .A2(_2292_),
    .B(_2297_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5337_ (.I(_2085_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5338_ (.A1(_2298_),
    .A2(_2089_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5339_ (.A1(_2097_),
    .A2(_2269_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5340_ (.A1(_2299_),
    .A2(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5341_ (.I(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_2302_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_2301_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5344_ (.I(_2304_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5345_ (.A1(\mod.registers.r4[0] ),
    .A2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5346_ (.A1(_2116_),
    .A2(_2303_),
    .B(_2306_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(\mod.registers.r4[1] ),
    .A2(_2305_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5348_ (.A1(_2127_),
    .A2(_2303_),
    .B(_2307_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5349_ (.A1(\mod.registers.r4[2] ),
    .A2(_2305_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5350_ (.A1(_2133_),
    .A2(_2303_),
    .B(_2308_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(\mod.registers.r4[3] ),
    .A2(_2305_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_2138_),
    .A2(_2303_),
    .B(_2309_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_2302_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5354_ (.I(_2304_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5355_ (.A1(\mod.registers.r4[4] ),
    .A2(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5356_ (.A1(_2145_),
    .A2(_2310_),
    .B(_2312_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5357_ (.A1(\mod.registers.r4[5] ),
    .A2(_2311_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5358_ (.A1(_2157_),
    .A2(_2310_),
    .B(_2313_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5359_ (.A1(\mod.registers.r4[6] ),
    .A2(_2311_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5360_ (.A1(_2167_),
    .A2(_2310_),
    .B(_2314_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(\mod.registers.r4[7] ),
    .A2(_2311_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5362_ (.A1(_2174_),
    .A2(_2310_),
    .B(_2315_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5363_ (.I(_2302_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_2304_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(\mod.registers.r4[8] ),
    .A2(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5366_ (.A1(_2184_),
    .A2(_2316_),
    .B(_2318_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5367_ (.A1(\mod.registers.r4[9] ),
    .A2(_2317_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5368_ (.A1(_2194_),
    .A2(_2316_),
    .B(_2319_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5369_ (.A1(\mod.registers.r4[10] ),
    .A2(_2317_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5370_ (.A1(_2202_),
    .A2(_2316_),
    .B(_2320_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5371_ (.A1(\mod.registers.r4[11] ),
    .A2(_2317_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5372_ (.A1(_2209_),
    .A2(_2316_),
    .B(_2321_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_2302_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5374_ (.I(_2304_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5375_ (.A1(\mod.registers.r4[12] ),
    .A2(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5376_ (.A1(_2217_),
    .A2(_2322_),
    .B(_2324_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5377_ (.A1(\mod.registers.r4[13] ),
    .A2(_2323_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5378_ (.A1(_2225_),
    .A2(_2322_),
    .B(_2325_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5379_ (.A1(\mod.registers.r4[14] ),
    .A2(_2323_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5380_ (.A1(_2231_),
    .A2(_2322_),
    .B(_2326_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5381_ (.A1(\mod.registers.r4[15] ),
    .A2(_2323_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5382_ (.A1(_2237_),
    .A2(_2322_),
    .B(_2327_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5383_ (.I(_2115_),
    .Z(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5384_ (.I(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5385_ (.A1(_2100_),
    .A2(_2299_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5386_ (.I(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5387_ (.I(_2331_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5388_ (.I(_2330_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5389_ (.I(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5390_ (.A1(\mod.registers.r5[0] ),
    .A2(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5391_ (.A1(_2329_),
    .A2(_2332_),
    .B(_2335_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5392_ (.I(_2126_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5393_ (.I(_2336_),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5394_ (.A1(\mod.registers.r5[1] ),
    .A2(_2334_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5395_ (.A1(_2337_),
    .A2(_2332_),
    .B(_2338_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5396_ (.I(_2132_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5397_ (.I(_2339_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5398_ (.A1(\mod.registers.r5[2] ),
    .A2(_2334_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5399_ (.A1(_2340_),
    .A2(_2332_),
    .B(_2341_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_2137_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_2342_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(\mod.registers.r5[3] ),
    .A2(_2334_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5403_ (.A1(_2343_),
    .A2(_2332_),
    .B(_2344_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5404_ (.I(_2144_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5405_ (.I(_2345_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5406_ (.I(_2331_),
    .Z(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_2333_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5408_ (.A1(\mod.registers.r5[4] ),
    .A2(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5409_ (.A1(_2346_),
    .A2(_2347_),
    .B(_2349_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_2156_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_2350_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5412_ (.A1(\mod.registers.r5[5] ),
    .A2(_2348_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5413_ (.A1(_2351_),
    .A2(_2347_),
    .B(_2352_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5414_ (.I(_2166_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5415_ (.I(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(\mod.registers.r5[6] ),
    .A2(_2348_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5417_ (.A1(_2354_),
    .A2(_2347_),
    .B(_2355_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5418_ (.I(_2173_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5419_ (.I(_2356_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(\mod.registers.r5[7] ),
    .A2(_2348_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(_2357_),
    .A2(_2347_),
    .B(_2358_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5422_ (.I(_2183_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5423_ (.I(_2359_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(_2331_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5425_ (.I(_2333_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5426_ (.A1(\mod.registers.r5[8] ),
    .A2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5427_ (.A1(_2360_),
    .A2(_2361_),
    .B(_2363_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_2193_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5429_ (.I(_2364_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(\mod.registers.r5[9] ),
    .A2(_2362_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5431_ (.A1(_2365_),
    .A2(_2361_),
    .B(_2366_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_2201_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5433_ (.I(_2367_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5434_ (.A1(\mod.registers.r5[10] ),
    .A2(_2362_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5435_ (.A1(_2368_),
    .A2(_2361_),
    .B(_2369_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5436_ (.I(_2208_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5437_ (.I(_2370_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(\mod.registers.r5[11] ),
    .A2(_2362_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5439_ (.A1(_2371_),
    .A2(_2361_),
    .B(_2372_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5440_ (.I(_2216_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_2373_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5442_ (.I(_2331_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5443_ (.I(_2333_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5444_ (.A1(\mod.registers.r5[12] ),
    .A2(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5445_ (.A1(_2374_),
    .A2(_2375_),
    .B(_2377_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5446_ (.I(_2224_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5447_ (.I(_2378_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5448_ (.A1(\mod.registers.r5[13] ),
    .A2(_2376_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5449_ (.A1(_2379_),
    .A2(_2375_),
    .B(_2380_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5450_ (.I(_2230_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5451_ (.I(_2381_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5452_ (.A1(\mod.registers.r5[14] ),
    .A2(_2376_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5453_ (.A1(_2382_),
    .A2(_2375_),
    .B(_2383_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_2236_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5455_ (.I(_2384_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5456_ (.A1(\mod.registers.r5[15] ),
    .A2(_2376_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5457_ (.A1(_2385_),
    .A2(_2375_),
    .B(_2386_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5458_ (.A1(_2241_),
    .A2(_2299_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5460_ (.I(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5461_ (.I(_2387_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5462_ (.I(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5463_ (.A1(\mod.registers.r6[0] ),
    .A2(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5464_ (.A1(_2329_),
    .A2(_2389_),
    .B(_2392_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5465_ (.A1(\mod.registers.r6[1] ),
    .A2(_2391_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5466_ (.A1(_2337_),
    .A2(_2389_),
    .B(_2393_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5467_ (.A1(\mod.registers.r6[2] ),
    .A2(_2391_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5468_ (.A1(_2340_),
    .A2(_2389_),
    .B(_2394_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5469_ (.A1(\mod.registers.r6[3] ),
    .A2(_2391_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5470_ (.A1(_2343_),
    .A2(_2389_),
    .B(_2395_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(_2388_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5472_ (.I(_2390_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5473_ (.A1(\mod.registers.r6[4] ),
    .A2(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5474_ (.A1(_2346_),
    .A2(_2396_),
    .B(_2398_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5475_ (.A1(\mod.registers.r6[5] ),
    .A2(_2397_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5476_ (.A1(_2351_),
    .A2(_2396_),
    .B(_2399_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(\mod.registers.r6[6] ),
    .A2(_2397_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5478_ (.A1(_2354_),
    .A2(_2396_),
    .B(_2400_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5479_ (.A1(\mod.registers.r6[7] ),
    .A2(_2397_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5480_ (.A1(_2357_),
    .A2(_2396_),
    .B(_2401_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5481_ (.I(_2388_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5482_ (.I(_2390_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5483_ (.A1(\mod.registers.r6[8] ),
    .A2(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5484_ (.A1(_2360_),
    .A2(_2402_),
    .B(_2404_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5485_ (.A1(\mod.registers.r6[9] ),
    .A2(_2403_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5486_ (.A1(_2365_),
    .A2(_2402_),
    .B(_2405_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5487_ (.A1(\mod.registers.r6[10] ),
    .A2(_2403_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5488_ (.A1(_2368_),
    .A2(_2402_),
    .B(_2406_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(\mod.registers.r6[11] ),
    .A2(_2403_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5490_ (.A1(_2371_),
    .A2(_2402_),
    .B(_2407_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5491_ (.I(_2388_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5492_ (.I(_2390_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5493_ (.A1(\mod.registers.r6[12] ),
    .A2(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5494_ (.A1(_2374_),
    .A2(_2408_),
    .B(_2410_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5495_ (.A1(\mod.registers.r6[13] ),
    .A2(_2409_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5496_ (.A1(_2379_),
    .A2(_2408_),
    .B(_2411_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5497_ (.A1(\mod.registers.r6[14] ),
    .A2(_2409_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5498_ (.A1(_2382_),
    .A2(_2408_),
    .B(_2412_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5499_ (.A1(\mod.registers.r6[15] ),
    .A2(_2409_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5500_ (.A1(_2385_),
    .A2(_2408_),
    .B(_2413_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5501_ (.A1(_2270_),
    .A2(_2299_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5502_ (.I(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5503_ (.I(_2415_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5504_ (.I(_2414_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5505_ (.I(_2417_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5506_ (.A1(\mod.registers.r7[0] ),
    .A2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5507_ (.A1(_2329_),
    .A2(_2416_),
    .B(_2419_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5508_ (.A1(\mod.registers.r7[1] ),
    .A2(_2418_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5509_ (.A1(_2337_),
    .A2(_2416_),
    .B(_2420_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(\mod.registers.r7[2] ),
    .A2(_2418_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5511_ (.A1(_2340_),
    .A2(_2416_),
    .B(_2421_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(\mod.registers.r7[3] ),
    .A2(_2418_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5513_ (.A1(_2343_),
    .A2(_2416_),
    .B(_2422_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5514_ (.I(_2415_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5515_ (.I(_2417_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5516_ (.A1(\mod.registers.r7[4] ),
    .A2(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5517_ (.A1(_2346_),
    .A2(_2423_),
    .B(_2425_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5518_ (.A1(\mod.registers.r7[5] ),
    .A2(_2424_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5519_ (.A1(_2351_),
    .A2(_2423_),
    .B(_2426_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(\mod.registers.r7[6] ),
    .A2(_2424_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_2354_),
    .A2(_2423_),
    .B(_2427_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5522_ (.A1(\mod.registers.r7[7] ),
    .A2(_2424_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5523_ (.A1(_2357_),
    .A2(_2423_),
    .B(_2428_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5524_ (.I(_2415_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5525_ (.I(_2417_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5526_ (.A1(\mod.registers.r7[8] ),
    .A2(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5527_ (.A1(_2360_),
    .A2(_2429_),
    .B(_2431_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5528_ (.A1(\mod.registers.r7[9] ),
    .A2(_2430_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5529_ (.A1(_2365_),
    .A2(_2429_),
    .B(_2432_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5530_ (.A1(\mod.registers.r7[10] ),
    .A2(_2430_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5531_ (.A1(_2368_),
    .A2(_2429_),
    .B(_2433_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5532_ (.A1(\mod.registers.r7[11] ),
    .A2(_2430_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5533_ (.A1(_2371_),
    .A2(_2429_),
    .B(_2434_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5534_ (.I(_2415_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5535_ (.I(_2417_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5536_ (.A1(\mod.registers.r7[12] ),
    .A2(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5537_ (.A1(_2374_),
    .A2(_2435_),
    .B(_2437_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5538_ (.A1(\mod.registers.r7[13] ),
    .A2(_2436_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5539_ (.A1(_2379_),
    .A2(_2435_),
    .B(_2438_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5540_ (.A1(\mod.registers.r7[14] ),
    .A2(_2436_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5541_ (.A1(_2382_),
    .A2(_2435_),
    .B(_2439_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5542_ (.A1(\mod.registers.r7[15] ),
    .A2(_2436_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5543_ (.A1(_2385_),
    .A2(_2435_),
    .B(_2440_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5544_ (.I(_2089_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5545_ (.A1(_2085_),
    .A2(_2441_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5546_ (.A1(_2300_),
    .A2(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5547_ (.I(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5548_ (.I(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5549_ (.I(_2443_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5550_ (.I(_2446_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(\mod.registers.r8[0] ),
    .A2(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5552_ (.A1(_2329_),
    .A2(_2445_),
    .B(_2448_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5553_ (.A1(\mod.registers.r8[1] ),
    .A2(_2447_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5554_ (.A1(_2337_),
    .A2(_2445_),
    .B(_2449_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5555_ (.A1(\mod.registers.r8[2] ),
    .A2(_2447_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5556_ (.A1(_2340_),
    .A2(_2445_),
    .B(_2450_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5557_ (.A1(\mod.registers.r8[3] ),
    .A2(_2447_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5558_ (.A1(_2343_),
    .A2(_2445_),
    .B(_2451_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5559_ (.I(_2444_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5560_ (.I(_2446_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5561_ (.A1(\mod.registers.r8[4] ),
    .A2(_2453_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5562_ (.A1(_2346_),
    .A2(_2452_),
    .B(_2454_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5563_ (.A1(\mod.registers.r8[5] ),
    .A2(_2453_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5564_ (.A1(_2351_),
    .A2(_2452_),
    .B(_2455_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5565_ (.A1(\mod.registers.r8[6] ),
    .A2(_2453_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5566_ (.A1(_2354_),
    .A2(_2452_),
    .B(_2456_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5567_ (.A1(\mod.registers.r8[7] ),
    .A2(_2453_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5568_ (.A1(_2357_),
    .A2(_2452_),
    .B(_2457_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_2444_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5570_ (.I(_2446_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5571_ (.A1(\mod.registers.r8[8] ),
    .A2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5572_ (.A1(_2360_),
    .A2(_2458_),
    .B(_2460_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5573_ (.A1(\mod.registers.r8[9] ),
    .A2(_2459_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5574_ (.A1(_2365_),
    .A2(_2458_),
    .B(_2461_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5575_ (.A1(\mod.registers.r8[10] ),
    .A2(_2459_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5576_ (.A1(_2368_),
    .A2(_2458_),
    .B(_2462_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5577_ (.A1(\mod.registers.r8[11] ),
    .A2(_2459_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5578_ (.A1(_2371_),
    .A2(_2458_),
    .B(_2463_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_2444_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5580_ (.I(_2446_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5581_ (.A1(\mod.registers.r8[12] ),
    .A2(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5582_ (.A1(_2374_),
    .A2(_2464_),
    .B(_2466_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5583_ (.A1(\mod.registers.r8[13] ),
    .A2(_2465_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5584_ (.A1(_2379_),
    .A2(_2464_),
    .B(_2467_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5585_ (.A1(\mod.registers.r8[14] ),
    .A2(_2465_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5586_ (.A1(_2382_),
    .A2(_2464_),
    .B(_2468_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5587_ (.A1(\mod.registers.r8[15] ),
    .A2(_2465_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5588_ (.A1(_2385_),
    .A2(_2464_),
    .B(_2469_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5589_ (.I(_2115_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5590_ (.A1(_2100_),
    .A2(_2442_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5591_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5593_ (.I(_2471_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5594_ (.I(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5595_ (.A1(\mod.registers.r9[0] ),
    .A2(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5596_ (.A1(_2470_),
    .A2(_2473_),
    .B(_2476_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5597_ (.I(_2126_),
    .Z(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(\mod.registers.r9[1] ),
    .A2(_2475_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5599_ (.A1(_2477_),
    .A2(_2473_),
    .B(_2478_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5600_ (.I(_2132_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5601_ (.A1(\mod.registers.r9[2] ),
    .A2(_2475_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5602_ (.A1(_2479_),
    .A2(_2473_),
    .B(_2480_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5603_ (.I(_2137_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5604_ (.A1(\mod.registers.r9[3] ),
    .A2(_2475_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5605_ (.A1(_2481_),
    .A2(_2473_),
    .B(_2482_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_2144_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5607_ (.I(_2472_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5608_ (.I(_2474_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5609_ (.A1(\mod.registers.r9[4] ),
    .A2(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5610_ (.A1(_2483_),
    .A2(_2484_),
    .B(_2486_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(_2156_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5612_ (.A1(\mod.registers.r9[5] ),
    .A2(_2485_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5613_ (.A1(_2487_),
    .A2(_2484_),
    .B(_2488_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_2166_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5615_ (.A1(\mod.registers.r9[6] ),
    .A2(_2485_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5616_ (.A1(_2489_),
    .A2(_2484_),
    .B(_2490_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(_2173_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5618_ (.A1(\mod.registers.r9[7] ),
    .A2(_2485_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5619_ (.A1(_2491_),
    .A2(_2484_),
    .B(_2492_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5620_ (.I(_2183_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5621_ (.I(_2472_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5622_ (.I(_2474_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5623_ (.A1(\mod.registers.r9[8] ),
    .A2(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5624_ (.A1(_2493_),
    .A2(_2494_),
    .B(_2496_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(_2193_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5626_ (.A1(\mod.registers.r9[9] ),
    .A2(_2495_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5627_ (.A1(_2497_),
    .A2(_2494_),
    .B(_2498_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5628_ (.I(_2201_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5629_ (.A1(\mod.registers.r9[10] ),
    .A2(_2495_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5630_ (.A1(_2499_),
    .A2(_2494_),
    .B(_2500_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5631_ (.I(_2208_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5632_ (.A1(\mod.registers.r9[11] ),
    .A2(_2495_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5633_ (.A1(_2501_),
    .A2(_2494_),
    .B(_2502_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5634_ (.I(_2216_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5635_ (.I(_2472_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5636_ (.I(_2474_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5637_ (.A1(\mod.registers.r9[12] ),
    .A2(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5638_ (.A1(_2503_),
    .A2(_2504_),
    .B(_2506_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5639_ (.I(_2224_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5640_ (.A1(\mod.registers.r9[13] ),
    .A2(_2505_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5641_ (.A1(_2507_),
    .A2(_2504_),
    .B(_2508_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5642_ (.I(_2230_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5643_ (.A1(\mod.registers.r9[14] ),
    .A2(_2505_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_2509_),
    .A2(_2504_),
    .B(_2510_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5645_ (.I(_2236_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5646_ (.A1(\mod.registers.r9[15] ),
    .A2(_2505_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5647_ (.A1(_2511_),
    .A2(_2504_),
    .B(_2512_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5648_ (.A1(_2241_),
    .A2(_2442_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5649_ (.I(_2513_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5650_ (.I(_2514_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5651_ (.I(_2513_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5652_ (.I(_2516_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5653_ (.A1(\mod.registers.r10[0] ),
    .A2(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5654_ (.A1(_2470_),
    .A2(_2515_),
    .B(_2518_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(\mod.registers.r10[1] ),
    .A2(_2517_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5656_ (.A1(_2477_),
    .A2(_2515_),
    .B(_2519_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\mod.registers.r10[2] ),
    .A2(_2517_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_2479_),
    .A2(_2515_),
    .B(_2520_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5659_ (.A1(\mod.registers.r10[3] ),
    .A2(_2517_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5660_ (.A1(_2481_),
    .A2(_2515_),
    .B(_2521_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5661_ (.I(_2514_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5662_ (.I(_2516_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(\mod.registers.r10[4] ),
    .A2(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5664_ (.A1(_2483_),
    .A2(_2522_),
    .B(_2524_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5665_ (.A1(\mod.registers.r10[5] ),
    .A2(_2523_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5666_ (.A1(_2487_),
    .A2(_2522_),
    .B(_2525_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5667_ (.A1(\mod.registers.r10[6] ),
    .A2(_2523_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5668_ (.A1(_2489_),
    .A2(_2522_),
    .B(_2526_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5669_ (.A1(\mod.registers.r10[7] ),
    .A2(_2523_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5670_ (.A1(_2491_),
    .A2(_2522_),
    .B(_2527_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(_2514_),
    .Z(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5672_ (.I(_2516_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5673_ (.A1(\mod.registers.r10[8] ),
    .A2(_2529_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5674_ (.A1(_2493_),
    .A2(_2528_),
    .B(_2530_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5675_ (.A1(\mod.registers.r10[9] ),
    .A2(_2529_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5676_ (.A1(_2497_),
    .A2(_2528_),
    .B(_2531_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5677_ (.A1(\mod.registers.r10[10] ),
    .A2(_2529_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5678_ (.A1(_2499_),
    .A2(_2528_),
    .B(_2532_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5679_ (.A1(\mod.registers.r10[11] ),
    .A2(_2529_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5680_ (.A1(_2501_),
    .A2(_2528_),
    .B(_2533_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5681_ (.I(_2514_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_2516_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5683_ (.A1(\mod.registers.r10[12] ),
    .A2(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5684_ (.A1(_2503_),
    .A2(_2534_),
    .B(_2536_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5685_ (.A1(\mod.registers.r10[13] ),
    .A2(_2535_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5686_ (.A1(_2507_),
    .A2(_2534_),
    .B(_2537_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5687_ (.A1(\mod.registers.r10[14] ),
    .A2(_2535_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5688_ (.A1(_2509_),
    .A2(_2534_),
    .B(_2538_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5689_ (.A1(\mod.registers.r10[15] ),
    .A2(_2535_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5690_ (.A1(_2511_),
    .A2(_2534_),
    .B(_2539_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5691_ (.A1(_2270_),
    .A2(_2442_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5692_ (.I(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5693_ (.I(_2541_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_2540_),
    .Z(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_2543_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5696_ (.A1(\mod.registers.r11[0] ),
    .A2(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5697_ (.A1(_2470_),
    .A2(_2542_),
    .B(_2545_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5698_ (.A1(\mod.registers.r11[1] ),
    .A2(_2544_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_2477_),
    .A2(_2542_),
    .B(_2546_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5700_ (.A1(\mod.registers.r11[2] ),
    .A2(_2544_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5701_ (.A1(_2479_),
    .A2(_2542_),
    .B(_2547_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5702_ (.A1(\mod.registers.r11[3] ),
    .A2(_2544_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5703_ (.A1(_2481_),
    .A2(_2542_),
    .B(_2548_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5704_ (.I(_2541_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5705_ (.I(_2543_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5706_ (.A1(\mod.registers.r11[4] ),
    .A2(_2550_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5707_ (.A1(_2483_),
    .A2(_2549_),
    .B(_2551_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5708_ (.A1(\mod.registers.r11[5] ),
    .A2(_2550_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5709_ (.A1(_2487_),
    .A2(_2549_),
    .B(_2552_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(\mod.registers.r11[6] ),
    .A2(_2550_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5711_ (.A1(_2489_),
    .A2(_2549_),
    .B(_2553_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(\mod.registers.r11[7] ),
    .A2(_2550_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5713_ (.A1(_2491_),
    .A2(_2549_),
    .B(_2554_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5714_ (.I(_2541_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_2543_),
    .Z(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5716_ (.A1(\mod.registers.r11[8] ),
    .A2(_2556_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5717_ (.A1(_2493_),
    .A2(_2555_),
    .B(_2557_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(\mod.registers.r11[9] ),
    .A2(_2556_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5719_ (.A1(_2497_),
    .A2(_2555_),
    .B(_2558_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5720_ (.A1(\mod.registers.r11[10] ),
    .A2(_2556_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5721_ (.A1(_2499_),
    .A2(_2555_),
    .B(_2559_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5722_ (.A1(\mod.registers.r11[11] ),
    .A2(_2556_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5723_ (.A1(_2501_),
    .A2(_2555_),
    .B(_2560_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5724_ (.I(_2541_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5725_ (.I(_2543_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5726_ (.A1(\mod.registers.r11[12] ),
    .A2(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5727_ (.A1(_2503_),
    .A2(_2561_),
    .B(_2563_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5728_ (.A1(\mod.registers.r11[13] ),
    .A2(_2562_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5729_ (.A1(_2507_),
    .A2(_2561_),
    .B(_2564_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(\mod.registers.r11[14] ),
    .A2(_2562_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5731_ (.A1(_2509_),
    .A2(_2561_),
    .B(_2565_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5732_ (.A1(\mod.registers.r11[15] ),
    .A2(_2562_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5733_ (.A1(_2511_),
    .A2(_2561_),
    .B(_2566_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5734_ (.A1(_2298_),
    .A2(_2441_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5735_ (.A1(_2300_),
    .A2(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5736_ (.I(_2568_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_2569_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5738_ (.I(_2568_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5739_ (.I(_2571_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5740_ (.A1(\mod.registers.r12[0] ),
    .A2(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5741_ (.A1(_2470_),
    .A2(_2570_),
    .B(_2573_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5742_ (.A1(\mod.registers.r12[1] ),
    .A2(_2572_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5743_ (.A1(_2477_),
    .A2(_2570_),
    .B(_2574_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(\mod.registers.r12[2] ),
    .A2(_2572_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5745_ (.A1(_2479_),
    .A2(_2570_),
    .B(_2575_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5746_ (.A1(\mod.registers.r12[3] ),
    .A2(_2572_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5747_ (.A1(_2481_),
    .A2(_2570_),
    .B(_2576_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5748_ (.I(_2569_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_2571_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5750_ (.A1(\mod.registers.r12[4] ),
    .A2(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5751_ (.A1(_2483_),
    .A2(_2577_),
    .B(_2579_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5752_ (.A1(\mod.registers.r12[5] ),
    .A2(_2578_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5753_ (.A1(_2487_),
    .A2(_2577_),
    .B(_2580_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5754_ (.A1(\mod.registers.r12[6] ),
    .A2(_2578_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5755_ (.A1(_2489_),
    .A2(_2577_),
    .B(_2581_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(\mod.registers.r12[7] ),
    .A2(_2578_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5757_ (.A1(_2491_),
    .A2(_2577_),
    .B(_2582_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5758_ (.I(_2569_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5759_ (.I(_2571_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(\mod.registers.r12[8] ),
    .A2(_2584_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5761_ (.A1(_2493_),
    .A2(_2583_),
    .B(_2585_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5762_ (.A1(\mod.registers.r12[9] ),
    .A2(_2584_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5763_ (.A1(_2497_),
    .A2(_2583_),
    .B(_2586_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5764_ (.A1(\mod.registers.r12[10] ),
    .A2(_2584_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5765_ (.A1(_2499_),
    .A2(_2583_),
    .B(_2587_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(\mod.registers.r12[11] ),
    .A2(_2584_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5767_ (.A1(_2501_),
    .A2(_2583_),
    .B(_2588_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5768_ (.I(_2569_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5769_ (.I(_2571_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5770_ (.A1(\mod.registers.r12[12] ),
    .A2(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5771_ (.A1(_2503_),
    .A2(_2589_),
    .B(_2591_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5772_ (.A1(\mod.registers.r12[13] ),
    .A2(_2590_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5773_ (.A1(_2507_),
    .A2(_2589_),
    .B(_2592_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5774_ (.A1(\mod.registers.r12[14] ),
    .A2(_2590_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5775_ (.A1(_2509_),
    .A2(_2589_),
    .B(_2593_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5776_ (.A1(\mod.registers.r12[15] ),
    .A2(_2590_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5777_ (.A1(_2511_),
    .A2(_2589_),
    .B(_2594_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5778_ (.A1(_2100_),
    .A2(_2567_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5779_ (.I(_2595_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_2596_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5781_ (.I(_2595_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5782_ (.I(_2598_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5783_ (.A1(\mod.registers.r13[0] ),
    .A2(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5784_ (.A1(_2328_),
    .A2(_2597_),
    .B(_2600_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(\mod.registers.r13[1] ),
    .A2(_2599_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5786_ (.A1(_2336_),
    .A2(_2597_),
    .B(_2601_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(\mod.registers.r13[2] ),
    .A2(_2599_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5788_ (.A1(_2339_),
    .A2(_2597_),
    .B(_2602_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5789_ (.A1(\mod.registers.r13[3] ),
    .A2(_2599_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5790_ (.A1(_2342_),
    .A2(_2597_),
    .B(_2603_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5791_ (.I(_2596_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(_2598_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5793_ (.A1(\mod.registers.r13[4] ),
    .A2(_2605_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5794_ (.A1(_2345_),
    .A2(_2604_),
    .B(_2606_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5795_ (.A1(\mod.registers.r13[5] ),
    .A2(_2605_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5796_ (.A1(_2350_),
    .A2(_2604_),
    .B(_2607_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(\mod.registers.r13[6] ),
    .A2(_2605_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5798_ (.A1(_2353_),
    .A2(_2604_),
    .B(_2608_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5799_ (.A1(\mod.registers.r13[7] ),
    .A2(_2605_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5800_ (.A1(_2356_),
    .A2(_2604_),
    .B(_2609_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5801_ (.I(_2596_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5802_ (.I(_2598_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5803_ (.A1(\mod.registers.r13[8] ),
    .A2(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5804_ (.A1(_2359_),
    .A2(_2610_),
    .B(_2612_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5805_ (.A1(\mod.registers.r13[9] ),
    .A2(_2611_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5806_ (.A1(_2364_),
    .A2(_2610_),
    .B(_2613_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(\mod.registers.r13[10] ),
    .A2(_2611_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5808_ (.A1(_2367_),
    .A2(_2610_),
    .B(_2614_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5809_ (.A1(\mod.registers.r13[11] ),
    .A2(_2611_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5810_ (.A1(_2370_),
    .A2(_2610_),
    .B(_2615_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5811_ (.I(_2596_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5812_ (.I(_2598_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5813_ (.A1(\mod.registers.r13[12] ),
    .A2(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5814_ (.A1(_2373_),
    .A2(_2616_),
    .B(_2618_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(\mod.registers.r13[13] ),
    .A2(_2617_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5816_ (.A1(_2378_),
    .A2(_2616_),
    .B(_2619_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(\mod.registers.r13[14] ),
    .A2(_2617_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(_2381_),
    .A2(_2616_),
    .B(_2620_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5819_ (.A1(\mod.registers.r13[15] ),
    .A2(_2617_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5820_ (.A1(_2384_),
    .A2(_2616_),
    .B(_2621_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5821_ (.A1(_2241_),
    .A2(_2567_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5822_ (.I(_2622_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5823_ (.I(_2623_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5824_ (.I(_2622_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5825_ (.I(_2625_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5826_ (.A1(\mod.registers.r14[0] ),
    .A2(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5827_ (.A1(_2328_),
    .A2(_2624_),
    .B(_2627_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(\mod.registers.r14[1] ),
    .A2(_2626_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5829_ (.A1(_2336_),
    .A2(_2624_),
    .B(_2628_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5830_ (.A1(\mod.registers.r14[2] ),
    .A2(_2626_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5831_ (.A1(_2339_),
    .A2(_2624_),
    .B(_2629_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5832_ (.A1(\mod.registers.r14[3] ),
    .A2(_2626_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5833_ (.A1(_2342_),
    .A2(_2624_),
    .B(_2630_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5834_ (.I(_2623_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5835_ (.I(_2625_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5836_ (.A1(\mod.registers.r14[4] ),
    .A2(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5837_ (.A1(_2345_),
    .A2(_2631_),
    .B(_2633_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5838_ (.A1(\mod.registers.r14[5] ),
    .A2(_2632_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5839_ (.A1(_2350_),
    .A2(_2631_),
    .B(_2634_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(\mod.registers.r14[6] ),
    .A2(_2632_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5841_ (.A1(_2353_),
    .A2(_2631_),
    .B(_2635_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(\mod.registers.r14[7] ),
    .A2(_2632_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5843_ (.A1(_2356_),
    .A2(_2631_),
    .B(_2636_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_2623_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5845_ (.I(_2625_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(\mod.registers.r14[8] ),
    .A2(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5847_ (.A1(_2359_),
    .A2(_2637_),
    .B(_2639_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5848_ (.A1(\mod.registers.r14[9] ),
    .A2(_2638_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5849_ (.A1(_2364_),
    .A2(_2637_),
    .B(_2640_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5850_ (.A1(\mod.registers.r14[10] ),
    .A2(_2638_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5851_ (.A1(_2367_),
    .A2(_2637_),
    .B(_2641_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5852_ (.A1(\mod.registers.r14[11] ),
    .A2(_2638_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5853_ (.A1(_2370_),
    .A2(_2637_),
    .B(_2642_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5854_ (.I(_2623_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5855_ (.I(_2625_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5856_ (.A1(\mod.registers.r14[12] ),
    .A2(_2644_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5857_ (.A1(_2373_),
    .A2(_2643_),
    .B(_2645_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5858_ (.A1(\mod.registers.r14[13] ),
    .A2(_2644_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5859_ (.A1(_2378_),
    .A2(_2643_),
    .B(_2646_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5860_ (.A1(\mod.registers.r14[14] ),
    .A2(_2644_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5861_ (.A1(_2381_),
    .A2(_2643_),
    .B(_2647_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5862_ (.A1(\mod.registers.r14[15] ),
    .A2(_2644_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5863_ (.A1(_2384_),
    .A2(_2643_),
    .B(_2648_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5864_ (.I(net11),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5865_ (.I(_2649_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_2650_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5867_ (.I(_2651_),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5868_ (.I(_2652_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5869_ (.I(_2652_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5870_ (.I(_2652_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5871_ (.A1(_1890_),
    .A2(_1828_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5872_ (.A1(\mod.valid0 ),
    .A2(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5873_ (.I(net12),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5874_ (.A1(_2655_),
    .A2(_1828_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5875_ (.I(_2656_),
    .Z(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5876_ (.I(_2657_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5877_ (.I(_2649_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5878_ (.I(_2659_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5879_ (.A1(_2654_),
    .A2(_2658_),
    .B(_2660_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5880_ (.I(_2093_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5881_ (.A1(\mod.valid0 ),
    .A2(_2653_),
    .A3(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5882_ (.I(_2662_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5883_ (.I(_2663_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5884_ (.I(_2656_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5885_ (.A1(\mod.valid1 ),
    .A2(_2653_),
    .A3(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5886_ (.A1(_2664_),
    .A2(_2666_),
    .B(_2660_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5887_ (.I(_2655_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5888_ (.I(_2667_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_2668_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5890_ (.I(_2667_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5891_ (.I(_2080_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5892_ (.A1(_2670_),
    .A2(\mod.pc0[0] ),
    .B(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5893_ (.A1(_2669_),
    .A2(_1847_),
    .B(_2672_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5894_ (.I(_2080_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5895_ (.A1(_2670_),
    .A2(\mod.pc0[1] ),
    .B(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5896_ (.A1(_2669_),
    .A2(_1871_),
    .B(_2674_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5897_ (.I(_2667_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5898_ (.A1(_2675_),
    .A2(_1886_),
    .A3(_1894_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5899_ (.I(_2655_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5900_ (.I(_2677_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5901_ (.A1(_2678_),
    .A2(\mod.pc0[2] ),
    .B(_0003_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5902_ (.A1(_2676_),
    .A2(_2679_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5903_ (.A1(_2675_),
    .A2(_1908_),
    .A3(_1912_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5904_ (.A1(_2678_),
    .A2(\mod.pc0[3] ),
    .B(_0003_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5905_ (.A1(_2680_),
    .A2(_2681_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5906_ (.A1(_2675_),
    .A2(_1926_),
    .A3(_1930_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5907_ (.I(_2667_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_2080_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5909_ (.A1(_2683_),
    .A2(\mod.pc0[4] ),
    .B(_2684_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5910_ (.A1(_2682_),
    .A2(_2685_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5911_ (.A1(_2668_),
    .A2(\mod.pc0[5] ),
    .B(_2673_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5912_ (.A1(_2669_),
    .A2(_1947_),
    .B(_2686_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5913_ (.A1(_2675_),
    .A2(_1960_),
    .A3(_1964_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5914_ (.A1(_2683_),
    .A2(\mod.pc0[6] ),
    .B(_2684_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5915_ (.A1(_2687_),
    .A2(_2688_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5916_ (.I(_2677_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5917_ (.A1(_2689_),
    .A2(_1977_),
    .A3(_1980_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5918_ (.A1(_2683_),
    .A2(\mod.pc0[7] ),
    .B(_2684_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_2690_),
    .A2(_2691_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5920_ (.A1(_2668_),
    .A2(\mod.pc0[8] ),
    .B(_2673_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5921_ (.A1(_2669_),
    .A2(_1995_),
    .B(_2692_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5922_ (.A1(_2689_),
    .A2(_2013_),
    .A3(_2016_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5923_ (.A1(_2683_),
    .A2(\mod.pc0[9] ),
    .B(_2684_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5924_ (.A1(_2693_),
    .A2(_2694_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5925_ (.A1(_2668_),
    .A2(\mod.pc0[10] ),
    .B(_2673_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5926_ (.A1(_2678_),
    .A2(_2031_),
    .B(_2695_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5927_ (.A1(_2670_),
    .A2(\mod.pc0[11] ),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5928_ (.I(_2677_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5929_ (.A1(_2697_),
    .A2(_2045_),
    .B(_2671_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5930_ (.A1(_2696_),
    .A2(_2698_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5931_ (.A1(_2689_),
    .A2(_2054_),
    .A3(_2057_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5932_ (.A1(_2670_),
    .A2(\mod.pc0[12] ),
    .B(_2671_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5933_ (.A1(_2699_),
    .A2(_2700_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5934_ (.A1(_2689_),
    .A2(_2068_),
    .A3(_2071_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5935_ (.A1(\mod.pc0[13] ),
    .A2(_2678_),
    .B(_2671_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5936_ (.A1(_2701_),
    .A2(_2702_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5937_ (.I(\mod.pc[0] ),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5938_ (.A1(_1868_),
    .A2(_1928_),
    .B(_2655_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5939_ (.I(_2704_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_2705_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5941_ (.I(_2704_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5942_ (.A1(_1739_),
    .A2(_1840_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5943_ (.I(_2079_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5944_ (.I(_2709_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5945_ (.I(_2710_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5946_ (.A1(_2707_),
    .A2(_2708_),
    .B(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5947_ (.A1(_2703_),
    .A2(_2706_),
    .B(_2712_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5948_ (.A1(_2697_),
    .A2(_1961_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5949_ (.I(_2713_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5950_ (.A1(_1855_),
    .A2(_1829_),
    .A3(_1866_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5951_ (.A1(_1869_),
    .A2(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5952_ (.A1(_2708_),
    .A2(_2716_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5953_ (.A1(\mod.pc[1] ),
    .A2(_2714_),
    .B(_2711_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5954_ (.A1(_2714_),
    .A2(_2717_),
    .B(_2718_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5955_ (.I(_2705_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5956_ (.I(\mod.pc[1] ),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5957_ (.A1(_2720_),
    .A2(_1856_),
    .B1(_1739_),
    .B2(_1840_),
    .C(_2715_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5958_ (.I(_2721_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5959_ (.A1(_1837_),
    .A2(_1839_),
    .B(\mod.pc[2] ),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5960_ (.A1(_1886_),
    .A2(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5961_ (.A1(_2722_),
    .A2(_2724_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5962_ (.A1(_2705_),
    .A2(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5963_ (.I(_2650_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5964_ (.A1(_1888_),
    .A2(_2719_),
    .B(_2726_),
    .C(_2727_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5965_ (.I(\mod.pc[3] ),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5966_ (.A1(_1886_),
    .A2(_2723_),
    .B1(_1908_),
    .B2(_1910_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5967_ (.A1(_2722_),
    .A2(_2729_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5968_ (.A1(_1908_),
    .A2(_1910_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5969_ (.A1(_2722_),
    .A2(_2724_),
    .B(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5970_ (.A1(_2730_),
    .A2(_2732_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5971_ (.A1(_2707_),
    .A2(_2733_),
    .B(_2711_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5972_ (.A1(_2728_),
    .A2(_2706_),
    .B(_2734_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5973_ (.A1(_1942_),
    .A2(_1943_),
    .B(\mod.pc[4] ),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5974_ (.A1(_1926_),
    .A2(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5975_ (.A1(_2721_),
    .A2(_2729_),
    .A3(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5976_ (.A1(_2730_),
    .A2(_2736_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5977_ (.I(_2704_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5978_ (.A1(_2737_),
    .A2(_2738_),
    .B(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(_2650_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5980_ (.A1(_1927_),
    .A2(_2719_),
    .B(_2740_),
    .C(_2741_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5981_ (.I(\mod.pc[5] ),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(_1941_),
    .A2(_1944_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5983_ (.A1(_2737_),
    .A2(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5984_ (.A1(_2707_),
    .A2(_2744_),
    .B(_2711_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5985_ (.A1(_2742_),
    .A2(_2706_),
    .B(_2745_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5986_ (.I(\mod.pc[6] ),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5987_ (.A1(_1926_),
    .A2(_2735_),
    .B1(_1941_),
    .B2(_1944_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5988_ (.A1(_2722_),
    .A2(_2729_),
    .A3(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5989_ (.A1(_1960_),
    .A2(_1962_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5990_ (.A1(_2748_),
    .A2(_2749_),
    .Z(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5991_ (.I(_2710_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5992_ (.A1(_2707_),
    .A2(_2750_),
    .B(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5993_ (.A1(_2746_),
    .A2(_2706_),
    .B(_2752_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5994_ (.I(\mod.pc[7] ),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5995_ (.A1(_2748_),
    .A2(_2749_),
    .B(_1977_),
    .C(_1978_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5996_ (.A1(_1960_),
    .A2(_1962_),
    .B1(_1977_),
    .B2(_1978_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5997_ (.A1(_2721_),
    .A2(_2729_),
    .A3(_2747_),
    .A4(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_2756_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5999_ (.A1(_2754_),
    .A2(_2757_),
    .B(_2739_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6000_ (.A1(_2753_),
    .A2(_2719_),
    .B(_2758_),
    .C(_2741_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(\mod.pc[8] ),
    .A2(_1857_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6002_ (.A1(_2759_),
    .A2(_1994_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6003_ (.A1(_2756_),
    .A2(_2760_),
    .Z(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6004_ (.A1(_2705_),
    .A2(_2761_),
    .B(_2751_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6005_ (.A1(_1982_),
    .A2(_2719_),
    .B(_2762_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6006_ (.I(_2704_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6007_ (.A1(\mod.pc[9] ),
    .A2(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6008_ (.A1(_2757_),
    .A2(_2760_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6009_ (.I0(\mod.pc[9] ),
    .I1(_2012_),
    .S(_1842_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6010_ (.I0(\mod.pc[8] ),
    .I1(_1993_),
    .S(_1890_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6011_ (.A1(_2767_),
    .A2(_2766_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6012_ (.A1(_2765_),
    .A2(_2766_),
    .B1(_2768_),
    .B2(_2757_),
    .C(_2713_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6013_ (.A1(_2764_),
    .A2(_2769_),
    .B(_2660_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(\mod.pc[10] ),
    .A2(_2763_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(_2756_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6016_ (.A1(_2771_),
    .A2(_2768_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6017_ (.I0(\mod.pc[10] ),
    .I1(_2030_),
    .S(_1890_),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6018_ (.A1(_2767_),
    .A2(_2766_),
    .A3(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6019_ (.I(_2774_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6020_ (.A1(_2772_),
    .A2(_2773_),
    .B1(_2775_),
    .B2(_2757_),
    .C(_2713_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6021_ (.A1(_2770_),
    .A2(_2776_),
    .B(_2660_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6022_ (.I(\mod.pc[11] ),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6023_ (.A1(_2777_),
    .A2(_1891_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6024_ (.A1(_1891_),
    .A2(_2044_),
    .B(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6025_ (.A1(_2771_),
    .A2(_2775_),
    .A3(_2779_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6026_ (.A1(_2771_),
    .A2(_2775_),
    .B(_2779_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6027_ (.A1(_2780_),
    .A2(_2781_),
    .B(_2739_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6028_ (.A1(_2777_),
    .A2(_2763_),
    .B(_2782_),
    .C(_2741_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6029_ (.A1(_2756_),
    .A2(_2774_),
    .A3(_2779_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6030_ (.A1(\mod.pc[12] ),
    .A2(_1857_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6031_ (.A1(_2054_),
    .A2(_2784_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6032_ (.A1(_2783_),
    .A2(_2785_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6033_ (.A1(\mod.pc[12] ),
    .A2(_2714_),
    .B(_2751_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6034_ (.A1(_2714_),
    .A2(_2786_),
    .B(_2787_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6035_ (.A1(_2771_),
    .A2(_2775_),
    .A3(_2779_),
    .A4(_2785_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6036_ (.I(_2068_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6037_ (.A1(_2789_),
    .A2(_2070_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6038_ (.A1(_2788_),
    .A2(_2790_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6039_ (.A1(_2788_),
    .A2(_2790_),
    .B(_2739_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6040_ (.A1(_2069_),
    .A2(_2763_),
    .B1(_2791_),
    .B2(_2792_),
    .C(_2741_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6041_ (.I(_2661_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6042_ (.I(_2793_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6043_ (.I(_2794_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6044_ (.I(_2793_),
    .Z(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6045_ (.I(_2796_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6046_ (.A1(\mod.pc_1[0] ),
    .A2(_2797_),
    .B(_2751_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6047_ (.A1(_2703_),
    .A2(_2795_),
    .B(_2798_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6048_ (.I(_2710_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6049_ (.A1(\mod.pc_1[1] ),
    .A2(_2797_),
    .B(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6050_ (.A1(_2720_),
    .A2(_2795_),
    .B(_2800_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6051_ (.A1(\mod.pc_1[2] ),
    .A2(_2797_),
    .B(_2799_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6052_ (.A1(_1888_),
    .A2(_2795_),
    .B(_2801_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6053_ (.A1(\mod.pc_1[3] ),
    .A2(_2797_),
    .B(_2799_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6054_ (.A1(_2728_),
    .A2(_2795_),
    .B(_2802_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6055_ (.I(_2794_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6056_ (.I(_2793_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6057_ (.I(_2804_),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6058_ (.A1(\mod.pc_1[4] ),
    .A2(_2805_),
    .B(_2799_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6059_ (.A1(_1927_),
    .A2(_2803_),
    .B(_2806_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_2710_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6061_ (.A1(\mod.pc_1[5] ),
    .A2(_2805_),
    .B(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6062_ (.A1(_2742_),
    .A2(_2803_),
    .B(_2808_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6063_ (.A1(\mod.pc_1[6] ),
    .A2(_2805_),
    .B(_2807_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6064_ (.A1(_2746_),
    .A2(_2803_),
    .B(_2809_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6065_ (.A1(\mod.pc_1[7] ),
    .A2(_2805_),
    .B(_2807_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6066_ (.A1(_2753_),
    .A2(_2803_),
    .B(_2810_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6067_ (.I(_2794_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_2804_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6069_ (.A1(\mod.pc_1[8] ),
    .A2(_2812_),
    .B(_2807_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6070_ (.A1(_1982_),
    .A2(_2811_),
    .B(_2813_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6071_ (.I(_2709_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6072_ (.I(_2814_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6073_ (.A1(\mod.pc_1[9] ),
    .A2(_2812_),
    .B(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6074_ (.A1(_2014_),
    .A2(_2811_),
    .B(_2816_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6075_ (.A1(\mod.pc_1[10] ),
    .A2(_2812_),
    .B(_2815_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6076_ (.A1(_2019_),
    .A2(_2811_),
    .B(_2817_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6077_ (.A1(\mod.pc_1[11] ),
    .A2(_2812_),
    .B(_2815_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6078_ (.A1(_2777_),
    .A2(_2811_),
    .B(_2818_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6079_ (.I(_2794_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6080_ (.I(_2804_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6081_ (.A1(\mod.pc_1[12] ),
    .A2(_2820_),
    .B(_2815_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6082_ (.A1(_2055_),
    .A2(_2819_),
    .B(_2821_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6083_ (.I(_2814_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6084_ (.A1(\mod.pc_1[13] ),
    .A2(_2820_),
    .B(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6085_ (.A1(_2069_),
    .A2(_2819_),
    .B(_2823_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6086_ (.I(\mod.instr[0] ),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6087_ (.I(_2662_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6088_ (.I(_2825_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6089_ (.A1(\mod.des.des_dout[0] ),
    .A2(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6090_ (.I(net13),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(_2828_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6092_ (.I(_2649_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6093_ (.I(_2830_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6094_ (.A1(_2824_),
    .A2(_2664_),
    .B1(_2827_),
    .B2(_2829_),
    .C(_2831_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6095_ (.I(\mod.instr[1] ),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6096_ (.A1(\mod.des.des_dout[1] ),
    .A2(_2826_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6097_ (.A1(_2832_),
    .A2(_2664_),
    .B1(_2833_),
    .B2(_2829_),
    .C(_2831_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6098_ (.I(\mod.instr[2] ),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(_2825_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6100_ (.A1(\mod.des.des_dout[2] ),
    .A2(_2835_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6101_ (.A1(_2834_),
    .A2(_2664_),
    .B1(_2836_),
    .B2(_2829_),
    .C(_2831_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6102_ (.I(\mod.instr[3] ),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6103_ (.I(_2662_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6104_ (.I(_2838_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6105_ (.A1(\mod.des.des_dout[3] ),
    .A2(_2835_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6106_ (.A1(_2837_),
    .A2(_2839_),
    .B1(_2840_),
    .B2(_2829_),
    .C(_2831_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6107_ (.I(\mod.instr[4] ),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6108_ (.A1(\mod.des.des_dout[4] ),
    .A2(_2835_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_2828_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_2830_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6111_ (.A1(_2841_),
    .A2(_2839_),
    .B1(_2842_),
    .B2(_2843_),
    .C(_2844_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6112_ (.I(\mod.instr[5] ),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6113_ (.A1(\mod.des.des_dout[5] ),
    .A2(_2835_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6114_ (.A1(_2845_),
    .A2(_2839_),
    .B1(_2846_),
    .B2(_2843_),
    .C(_2844_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6115_ (.I(\mod.instr[6] ),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6116_ (.I(_2825_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6117_ (.A1(\mod.des.des_dout[6] ),
    .A2(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6118_ (.A1(_2847_),
    .A2(_2839_),
    .B1(_2849_),
    .B2(_2843_),
    .C(_2844_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6119_ (.I(\mod.instr[7] ),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6120_ (.I(_2663_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6121_ (.A1(\mod.des.des_dout[7] ),
    .A2(_2848_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6122_ (.A1(_2850_),
    .A2(_2851_),
    .B1(_2852_),
    .B2(_2843_),
    .C(_2844_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6123_ (.I(\mod.instr[8] ),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6124_ (.A1(\mod.des.des_dout[8] ),
    .A2(_2848_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6125_ (.I(_2828_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6126_ (.I(_2830_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6127_ (.A1(_2853_),
    .A2(_2851_),
    .B1(_2854_),
    .B2(_2855_),
    .C(_2856_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6128_ (.I(\mod.instr[9] ),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6129_ (.A1(\mod.des.des_dout[9] ),
    .A2(_2848_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6130_ (.A1(_2857_),
    .A2(_2851_),
    .B1(_2858_),
    .B2(_2855_),
    .C(_2856_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6131_ (.I(\mod.instr[10] ),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6132_ (.I(_2825_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6133_ (.A1(\mod.des.des_dout[10] ),
    .A2(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6134_ (.A1(_2859_),
    .A2(_2851_),
    .B1(_2861_),
    .B2(_2855_),
    .C(_2856_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6135_ (.I(\mod.instr[11] ),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6136_ (.I(_2663_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6137_ (.A1(\mod.des.des_dout[11] ),
    .A2(_2860_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6138_ (.A1(_2862_),
    .A2(_2863_),
    .B1(_2864_),
    .B2(_2855_),
    .C(_2856_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6139_ (.I(\mod.instr[12] ),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6140_ (.A1(\mod.des.des_dout[12] ),
    .A2(_2860_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6141_ (.I(net13),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_2830_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6143_ (.A1(_2865_),
    .A2(_2863_),
    .B1(_2866_),
    .B2(_2867_),
    .C(_2868_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6144_ (.I(\mod.instr[13] ),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6145_ (.A1(\mod.des.des_dout[13] ),
    .A2(_2860_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6146_ (.A1(_2869_),
    .A2(_2863_),
    .B1(_2870_),
    .B2(_2867_),
    .C(_2868_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6147_ (.I(\mod.instr[14] ),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6148_ (.I(_2662_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6149_ (.A1(\mod.des.des_dout[14] ),
    .A2(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6150_ (.A1(_2871_),
    .A2(_2863_),
    .B1(_2873_),
    .B2(_2867_),
    .C(_2868_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6151_ (.I(\mod.instr[15] ),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6152_ (.I(_2663_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6153_ (.A1(\mod.des.des_dout[15] ),
    .A2(_2872_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6154_ (.A1(_2874_),
    .A2(_2875_),
    .B1(_2876_),
    .B2(_2867_),
    .C(_2868_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6155_ (.I(\mod.instr[16] ),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6156_ (.A1(\mod.des.des_dout[16] ),
    .A2(_2872_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6157_ (.I(net13),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6158_ (.I(_2650_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6159_ (.A1(_2877_),
    .A2(_2875_),
    .B1(_2878_),
    .B2(_2879_),
    .C(_2880_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6160_ (.I(\mod.instr[17] ),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6161_ (.A1(\mod.des.des_dout[17] ),
    .A2(_2872_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6162_ (.A1(_2881_),
    .A2(_2875_),
    .B1(_2882_),
    .B2(_2879_),
    .C(_2880_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6163_ (.I(\mod.instr[18] ),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6164_ (.A1(\mod.des.des_dout[18] ),
    .A2(_2838_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6165_ (.A1(_2883_),
    .A2(_2875_),
    .B1(_2884_),
    .B2(_2879_),
    .C(_2880_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6166_ (.I(\mod.instr[19] ),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6167_ (.A1(\mod.des.des_dout[19] ),
    .A2(_2838_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6168_ (.A1(_2885_),
    .A2(_2826_),
    .B1(_2886_),
    .B2(_2879_),
    .C(_2880_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6169_ (.I(\mod.instr[20] ),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6170_ (.A1(\mod.des.des_dout[20] ),
    .A2(_2838_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6171_ (.I(_2649_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6172_ (.A1(_2887_),
    .A2(_2826_),
    .B1(_2888_),
    .B2(_2828_),
    .C(_2889_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6173_ (.A1(\mod.valid1 ),
    .A2(_2653_),
    .A3(_2661_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6174_ (.I(_2890_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6175_ (.I(_2656_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_2892_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6177_ (.A1(_2092_),
    .A2(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6178_ (.I(_2659_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6179_ (.A1(_2891_),
    .A2(_2894_),
    .B(_2895_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6180_ (.I(_2793_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6181_ (.I(_2896_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6182_ (.A1(_3114_),
    .A2(_2897_),
    .B1(_2891_),
    .B2(\mod.instr[0] ),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6183_ (.A1(_2652_),
    .A2(_2898_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_2889_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6185_ (.I(_2896_),
    .Z(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6186_ (.A1(_1860_),
    .A2(_2900_),
    .B1(_2891_),
    .B2(\mod.instr[1] ),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6187_ (.A1(_2899_),
    .A2(_2901_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6188_ (.A1(_3111_),
    .A2(_2900_),
    .B1(_2891_),
    .B2(\mod.instr[2] ),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6189_ (.A1(_2899_),
    .A2(_2902_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6190_ (.I(_2890_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6191_ (.I(_2903_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6192_ (.A1(\mod.instr_2[3] ),
    .A2(_2900_),
    .B1(_2904_),
    .B2(\mod.instr[3] ),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6193_ (.A1(_2899_),
    .A2(_2905_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6194_ (.A1(_1793_),
    .A2(_2900_),
    .B1(_2904_),
    .B2(\mod.instr[4] ),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6195_ (.A1(_2899_),
    .A2(_2906_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6196_ (.I(_2889_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6197_ (.I(_1804_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6198_ (.I(_2908_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6199_ (.I(_2896_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6200_ (.A1(_2909_),
    .A2(_2910_),
    .B1(_2904_),
    .B2(\mod.instr[5] ),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6201_ (.A1(_2907_),
    .A2(_2911_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6202_ (.A1(_1809_),
    .A2(_2910_),
    .B1(_2904_),
    .B2(\mod.instr[6] ),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6203_ (.A1(_2907_),
    .A2(_2912_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6204_ (.I(_2903_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6205_ (.A1(_1710_),
    .A2(_2910_),
    .B1(_2913_),
    .B2(\mod.instr[7] ),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6206_ (.A1(_2907_),
    .A2(_2914_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6207_ (.A1(_3119_),
    .A2(_2910_),
    .B1(_2913_),
    .B2(\mod.instr[8] ),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6208_ (.A1(_2907_),
    .A2(_2915_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6209_ (.I(_2889_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6210_ (.I(_2796_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6211_ (.A1(_1713_),
    .A2(_2917_),
    .B1(_2913_),
    .B2(\mod.instr[9] ),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6212_ (.A1(_2916_),
    .A2(_2918_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6213_ (.A1(_1749_),
    .A2(_2917_),
    .B1(_2913_),
    .B2(\mod.instr[10] ),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6214_ (.A1(_2916_),
    .A2(_2919_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6215_ (.I(_2890_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6216_ (.A1(_1750_),
    .A2(_2917_),
    .B1(_2920_),
    .B2(\mod.instr[11] ),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6217_ (.A1(_2916_),
    .A2(_2921_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6218_ (.A1(_0933_),
    .A2(_2917_),
    .B1(_2920_),
    .B2(\mod.instr[12] ),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6219_ (.A1(_2916_),
    .A2(_2922_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6220_ (.I(_2651_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_2796_),
    .Z(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6222_ (.A1(_0711_),
    .A2(_2924_),
    .B1(_2920_),
    .B2(\mod.instr[13] ),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6223_ (.A1(_2923_),
    .A2(_2925_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6224_ (.A1(_0695_),
    .A2(_2924_),
    .B1(_2920_),
    .B2(\mod.instr[14] ),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6225_ (.A1(_2923_),
    .A2(_2926_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6226_ (.I(_2890_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6227_ (.A1(_0501_),
    .A2(_2924_),
    .B1(_2927_),
    .B2(\mod.instr[15] ),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6228_ (.A1(_2923_),
    .A2(_2928_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6229_ (.A1(_0693_),
    .A2(_2924_),
    .B1(_2927_),
    .B2(\mod.instr[16] ),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6230_ (.A1(_2923_),
    .A2(_2929_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6231_ (.I(_2651_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_2796_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6233_ (.A1(_0657_),
    .A2(_2931_),
    .B1(_2927_),
    .B2(\mod.instr[17] ),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6234_ (.A1(_2930_),
    .A2(_2932_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6235_ (.A1(\mod.funct7[0] ),
    .A2(_2931_),
    .B1(_2927_),
    .B2(\mod.instr[18] ),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6236_ (.A1(_2930_),
    .A2(_2933_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6237_ (.A1(\mod.funct7[1] ),
    .A2(_2931_),
    .B1(_2903_),
    .B2(\mod.instr[19] ),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6238_ (.A1(_2930_),
    .A2(_2934_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6239_ (.A1(\mod.funct7[2] ),
    .A2(_2931_),
    .B1(_2903_),
    .B2(\mod.instr[20] ),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6240_ (.A1(_2930_),
    .A2(_2935_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6241_ (.I(_2892_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6242_ (.A1(\mod.pc_1[0] ),
    .A2(_2936_),
    .B(_2822_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6243_ (.A1(_1133_),
    .A2(_2658_),
    .B(_2937_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6244_ (.A1(\mod.pc_1[1] ),
    .A2(_2936_),
    .B(_2822_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6245_ (.A1(_0707_),
    .A2(_2658_),
    .B(_2938_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6246_ (.A1(\mod.pc_1[2] ),
    .A2(_2936_),
    .B(_2822_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6247_ (.A1(_0622_),
    .A2(_2658_),
    .B(_2939_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6248_ (.I(_2657_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6249_ (.I(_2892_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6250_ (.I(_2814_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6251_ (.A1(\mod.pc_1[3] ),
    .A2(_2941_),
    .B(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6252_ (.A1(_0676_),
    .A2(_2940_),
    .B(_2943_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6253_ (.A1(\mod.pc_1[4] ),
    .A2(_2941_),
    .B(_2942_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6254_ (.A1(_0568_),
    .A2(_2940_),
    .B(_2944_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6255_ (.A1(\mod.pc_1[5] ),
    .A2(_2941_),
    .B(_2942_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6256_ (.A1(_0591_),
    .A2(_2940_),
    .B(_2945_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6257_ (.A1(\mod.pc_1[6] ),
    .A2(_2941_),
    .B(_2942_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6258_ (.A1(_0453_),
    .A2(_2940_),
    .B(_2946_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6259_ (.I(_2657_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_2892_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_2814_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6262_ (.A1(\mod.pc_1[7] ),
    .A2(_2948_),
    .B(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6263_ (.A1(_0596_),
    .A2(_2947_),
    .B(_2950_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6264_ (.A1(\mod.pc_1[8] ),
    .A2(_2948_),
    .B(_2949_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6265_ (.A1(_0779_),
    .A2(_2947_),
    .B(_2951_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6266_ (.I(_2005_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6267_ (.A1(\mod.pc_1[9] ),
    .A2(_2948_),
    .B(_2949_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6268_ (.A1(_2952_),
    .A2(_2947_),
    .B(_2953_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6269_ (.A1(\mod.pc_1[10] ),
    .A2(_2948_),
    .B(_2949_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6270_ (.A1(_0911_),
    .A2(_2947_),
    .B(_2954_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(_2709_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6272_ (.A1(\mod.pc_1[11] ),
    .A2(_2665_),
    .B(_2955_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6273_ (.A1(_0878_),
    .A2(_2893_),
    .B(_2956_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6274_ (.A1(\mod.pc_1[12] ),
    .A2(_2665_),
    .B(_2955_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6275_ (.A1(_2062_),
    .A2(_2893_),
    .B(_2957_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6276_ (.A1(\mod.pc_1[13] ),
    .A2(_2665_),
    .B(_2955_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6277_ (.A1(_0957_),
    .A2(_2893_),
    .B(_2958_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6278_ (.A1(_2092_),
    .A2(_2896_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6279_ (.A1(\mod.valid_out3 ),
    .A2(_2091_),
    .A3(_2657_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6280_ (.A1(_2959_),
    .A2(_2960_),
    .B(_2895_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6281_ (.A1(net20),
    .A2(_2959_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6282_ (.I(_2804_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6283_ (.A1(_2092_),
    .A2(_1774_),
    .A3(_3123_),
    .A4(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6284_ (.A1(_2961_),
    .A2(_2963_),
    .B(_2895_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6285_ (.A1(\mod.ri_3 ),
    .A2(_2820_),
    .B(_2955_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6286_ (.A1(_0539_),
    .A2(_2819_),
    .B(_2964_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6287_ (.A1(_1774_),
    .A2(_2661_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6288_ (.A1(\mod.ins_ldr_3 ),
    .A2(_2936_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6289_ (.A1(_2965_),
    .A2(_2966_),
    .B(_2895_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6290_ (.I(_2709_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6291_ (.A1(\mod.rd_3[0] ),
    .A2(_2820_),
    .B(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6292_ (.A1(_1794_),
    .A2(_2819_),
    .B(_2968_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6293_ (.A1(\mod.rd_3[1] ),
    .A2(_2962_),
    .B(_2967_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6294_ (.A1(_1797_),
    .A2(_2897_),
    .B(_2969_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6295_ (.I(_0440_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6296_ (.A1(\mod.rd_3[2] ),
    .A2(_2962_),
    .B(_2967_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6297_ (.A1(_2970_),
    .A2(_2897_),
    .B(_2971_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6298_ (.A1(\mod.rd_3[3] ),
    .A2(_2962_),
    .B(_2967_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6299_ (.A1(_2086_),
    .A2(_2897_),
    .B(_2972_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6300_ (.A1(_2677_),
    .A2(_1744_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6302_ (.A1(_1753_),
    .A2(_0003_),
    .A3(_2974_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6303_ (.I(_2975_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(_1754_),
    .A2(_2974_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6305_ (.I(_1796_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6306_ (.A1(_1809_),
    .A2(_2965_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6307_ (.I(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6308_ (.A1(_2970_),
    .A2(_2977_),
    .A3(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6309_ (.I(_2659_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6310_ (.A1(_2976_),
    .A2(_2980_),
    .B(_2981_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6311_ (.A1(_1755_),
    .A2(_2974_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6312_ (.I(_1802_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6313_ (.A1(_2970_),
    .A2(_2983_),
    .A3(_2979_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6314_ (.A1(_2982_),
    .A2(_2984_),
    .B(_2981_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_1756_),
    .A2(_2974_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6316_ (.I(_1799_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6317_ (.A1(_2970_),
    .A2(_2986_),
    .A3(_2979_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6318_ (.A1(_2985_),
    .A2(_2987_),
    .B(_2981_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6319_ (.I(_2973_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6320_ (.A1(_1769_),
    .A2(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6321_ (.A1(_2909_),
    .A2(_1812_),
    .A3(_2979_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6322_ (.A1(_2989_),
    .A2(_2990_),
    .B(_2981_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6323_ (.A1(_1765_),
    .A2(_2988_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6324_ (.A1(_2909_),
    .A2(_2977_),
    .A3(_2978_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6325_ (.I(_2659_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6326_ (.A1(_2991_),
    .A2(_2992_),
    .B(_2993_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6327_ (.A1(_1768_),
    .A2(_2988_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6328_ (.A1(_2909_),
    .A2(_2983_),
    .A3(_2978_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6329_ (.A1(_2994_),
    .A2(_2995_),
    .B(_2993_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6330_ (.A1(_1767_),
    .A2(_2988_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6331_ (.I(_2908_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6332_ (.A1(_2997_),
    .A2(_2986_),
    .A3(_2978_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6333_ (.A1(_2996_),
    .A2(_2998_),
    .B(_2993_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6334_ (.I(_2651_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6335_ (.I(_2973_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6336_ (.A1(_2086_),
    .A2(_2908_),
    .A3(_2965_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6337_ (.A1(_1781_),
    .A2(_3000_),
    .B1(_3001_),
    .B2(_1812_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6338_ (.A1(_2999_),
    .A2(_3002_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6339_ (.A1(_1758_),
    .A2(_3000_),
    .B1(_3001_),
    .B2(_2977_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6340_ (.A1(_2999_),
    .A2(_3003_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6341_ (.A1(_1763_),
    .A2(_3000_),
    .B1(_3001_),
    .B2(_2983_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6342_ (.A1(_2999_),
    .A2(_3004_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6343_ (.A1(_1761_),
    .A2(_3000_),
    .B1(_3001_),
    .B2(_2986_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6344_ (.A1(_2999_),
    .A2(_3005_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6345_ (.I(_2973_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6346_ (.A1(_1745_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6347_ (.A1(_2086_),
    .A2(_2965_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6348_ (.A1(_2997_),
    .A2(_1812_),
    .A3(_3008_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6349_ (.A1(_3007_),
    .A2(_3009_),
    .B(_2993_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6350_ (.A1(_1746_),
    .A2(_3006_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6351_ (.A1(_2997_),
    .A2(_2977_),
    .A3(_3008_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6352_ (.A1(_3010_),
    .A2(_3011_),
    .B(_2727_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6353_ (.A1(_1747_),
    .A2(_3006_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6354_ (.A1(_2997_),
    .A2(_2983_),
    .A3(_3008_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6355_ (.A1(_3012_),
    .A2(_3013_),
    .B(_2727_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6356_ (.A1(_1748_),
    .A2(_3006_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6357_ (.A1(_2908_),
    .A2(_2986_),
    .A3(_3008_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6358_ (.A1(_3014_),
    .A2(_3015_),
    .B(_2727_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6359_ (.A1(_3092_),
    .A2(_3093_),
    .A3(\mod.des.des_counter[2] ),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6360_ (.I(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6361_ (.I0(\mod.des.des_dout[0] ),
    .I1(net16),
    .S(_3017_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6362_ (.I(_3018_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6363_ (.I0(\mod.des.des_dout[1] ),
    .I1(net17),
    .S(_3017_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_3019_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6365_ (.I0(\mod.des.des_dout[2] ),
    .I1(net18),
    .S(_3017_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6366_ (.I(_3020_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6367_ (.I0(\mod.des.des_dout[3] ),
    .I1(net19),
    .S(_3017_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6368_ (.I(_3021_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6369_ (.I(_3016_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6370_ (.I0(\mod.des.des_dout[4] ),
    .I1(net2),
    .S(_3022_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6371_ (.I(_3023_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6372_ (.I0(\mod.des.des_dout[5] ),
    .I1(net3),
    .S(_3022_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6373_ (.I(_3024_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6374_ (.I0(\mod.des.des_dout[6] ),
    .I1(net4),
    .S(_3022_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6375_ (.I(_3025_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6376_ (.I0(\mod.des.des_dout[7] ),
    .I1(net5),
    .S(_3022_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6377_ (.I(_3026_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6378_ (.I(_3016_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6379_ (.I0(\mod.des.des_dout[8] ),
    .I1(net6),
    .S(_3027_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6380_ (.I(_3028_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6381_ (.I0(\mod.des.des_dout[9] ),
    .I1(net7),
    .S(_3027_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6382_ (.I(_3029_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6383_ (.I0(\mod.des.des_dout[10] ),
    .I1(net8),
    .S(_3027_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6384_ (.I(_3030_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6385_ (.I0(\mod.des.des_dout[11] ),
    .I1(net9),
    .S(_3027_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6386_ (.I(_3031_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6387_ (.I0(\mod.des.des_dout[12] ),
    .I1(net10),
    .S(_3016_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6388_ (.I(_3032_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6389_ (.A1(_2270_),
    .A2(_2567_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6390_ (.I(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6391_ (.I(_3034_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6392_ (.I(_3033_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6393_ (.I(_3036_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6394_ (.A1(\mod.registers.r15[0] ),
    .A2(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6395_ (.A1(_2328_),
    .A2(_3035_),
    .B(_3038_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6396_ (.A1(\mod.registers.r15[1] ),
    .A2(_3037_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6397_ (.A1(_2336_),
    .A2(_3035_),
    .B(_3039_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6398_ (.A1(\mod.registers.r15[2] ),
    .A2(_3037_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6399_ (.A1(_2339_),
    .A2(_3035_),
    .B(_3040_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6400_ (.A1(\mod.registers.r15[3] ),
    .A2(_3037_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6401_ (.A1(_2342_),
    .A2(_3035_),
    .B(_3041_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6402_ (.I(_3034_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6403_ (.I(_3036_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6404_ (.A1(\mod.registers.r15[4] ),
    .A2(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6405_ (.A1(_2345_),
    .A2(_3042_),
    .B(_3044_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6406_ (.A1(\mod.registers.r15[5] ),
    .A2(_3043_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6407_ (.A1(_2350_),
    .A2(_3042_),
    .B(_3045_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6408_ (.A1(\mod.registers.r15[6] ),
    .A2(_3043_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6409_ (.A1(_2353_),
    .A2(_3042_),
    .B(_3046_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6410_ (.A1(\mod.registers.r15[7] ),
    .A2(_3043_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6411_ (.A1(_2356_),
    .A2(_3042_),
    .B(_3047_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6412_ (.I(_3034_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6413_ (.I(_3036_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6414_ (.A1(\mod.registers.r15[8] ),
    .A2(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6415_ (.A1(_2359_),
    .A2(_3048_),
    .B(_3050_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6416_ (.A1(\mod.registers.r15[9] ),
    .A2(_3049_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6417_ (.A1(_2364_),
    .A2(_3048_),
    .B(_3051_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6418_ (.A1(\mod.registers.r15[10] ),
    .A2(_3049_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6419_ (.A1(_2367_),
    .A2(_3048_),
    .B(_3052_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6420_ (.A1(\mod.registers.r15[11] ),
    .A2(_3049_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6421_ (.A1(_2370_),
    .A2(_3048_),
    .B(_3053_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_3034_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6423_ (.I(_3036_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6424_ (.A1(\mod.registers.r15[12] ),
    .A2(_3055_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6425_ (.A1(_2373_),
    .A2(_3054_),
    .B(_3056_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6426_ (.A1(\mod.registers.r15[13] ),
    .A2(_3055_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6427_ (.A1(_2378_),
    .A2(_3054_),
    .B(_3057_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(\mod.registers.r15[14] ),
    .A2(_3055_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6429_ (.A1(_2381_),
    .A2(_3054_),
    .B(_3058_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6430_ (.A1(\mod.registers.r15[15] ),
    .A2(_3055_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6431_ (.A1(_2384_),
    .A2(_3054_),
    .B(_3059_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6432_ (.A1(\mod.des.des_counter[2] ),
    .A2(_2074_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6433_ (.I(_3060_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6434_ (.I0(\mod.des.des_dout[13] ),
    .I1(net16),
    .S(_3061_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6435_ (.I(_3062_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6436_ (.I0(\mod.des.des_dout[14] ),
    .I1(net17),
    .S(_3061_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6437_ (.I(_3063_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6438_ (.I0(\mod.des.des_dout[15] ),
    .I1(net18),
    .S(_3061_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_3064_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6440_ (.I0(\mod.des.des_dout[16] ),
    .I1(net19),
    .S(_3061_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_3065_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6442_ (.I(_3060_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6443_ (.I0(\mod.des.des_dout[17] ),
    .I1(net2),
    .S(_3066_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_3067_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6445_ (.I0(\mod.des.des_dout[18] ),
    .I1(net3),
    .S(_3066_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6446_ (.I(_3068_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6447_ (.I0(\mod.des.des_dout[19] ),
    .I1(net4),
    .S(_3066_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6448_ (.I(_3069_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6449_ (.I0(\mod.des.des_dout[20] ),
    .I1(net5),
    .S(_3066_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6450_ (.I(_3070_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6451_ (.I(_3060_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6452_ (.I0(\mod.des.des_dout[21] ),
    .I1(net6),
    .S(_3071_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6453_ (.I(_3072_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6454_ (.I0(\mod.des.des_dout[22] ),
    .I1(net7),
    .S(_3071_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_3073_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6456_ (.I0(\mod.des.des_dout[23] ),
    .I1(net8),
    .S(_3071_),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6457_ (.I(_3074_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6458_ (.I0(\mod.des.des_dout[24] ),
    .I1(net9),
    .S(_3071_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6459_ (.I(_3075_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6460_ (.I0(\mod.des.des_dout[25] ),
    .I1(net10),
    .S(_3060_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6461_ (.I(_3076_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6462_ (.A1(\mod.des.des_counter[2] ),
    .A2(_2076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6463_ (.I(_3077_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6464_ (.I(_3078_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6465_ (.I0(\mod.des.des_dout[26] ),
    .I1(net16),
    .S(_3079_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6466_ (.I(_3080_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6467_ (.I0(\mod.des.des_dout[27] ),
    .I1(net17),
    .S(_3079_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6468_ (.I(_3081_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6469_ (.I0(\mod.des.des_dout[28] ),
    .I1(net18),
    .S(_3079_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6470_ (.I(_3082_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6471_ (.I0(\mod.des.des_dout[29] ),
    .I1(net19),
    .S(_3079_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6472_ (.I(_3083_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6473_ (.I(_3077_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6474_ (.I0(\mod.des.des_dout[30] ),
    .I1(net2),
    .S(_3084_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6475_ (.I(_3085_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6476_ (.I0(\mod.des.des_dout[31] ),
    .I1(net3),
    .S(_3084_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6477_ (.I(_3086_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6478_ (.I0(\mod.des.des_dout[32] ),
    .I1(net4),
    .S(_3084_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6479_ (.I(_3087_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6480_ (.I0(\mod.des.des_dout[33] ),
    .I1(net5),
    .S(_3084_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6481_ (.I(_3088_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6482_ (.I0(\mod.des.des_dout[34] ),
    .I1(net6),
    .S(_3078_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6483_ (.I(_3089_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6484_ (.I0(\mod.des.des_dout[35] ),
    .I1(net7),
    .S(_3078_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6485_ (.I(_3090_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6486_ (.I0(\mod.des.des_dout[36] ),
    .I1(net8),
    .S(_3078_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6487_ (.I(_3091_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6488_ (.D(_0121_),
    .RN(_0003_),
    .CLK(net201),
    .Q(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6489_ (.D(_0122_),
    .CLK(net116),
    .Q(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6490_ (.D(_0123_),
    .CLK(net118),
    .Q(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6491_ (.D(_0124_),
    .CLK(net115),
    .Q(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6492_ (.D(_0125_),
    .CLK(net117),
    .Q(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6493_ (.D(_0126_),
    .CLK(net100),
    .Q(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6494_ (.D(_0127_),
    .CLK(net98),
    .Q(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6495_ (.D(_0128_),
    .CLK(net100),
    .Q(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6496_ (.D(_0129_),
    .CLK(net99),
    .Q(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6497_ (.D(_0130_),
    .CLK(net43),
    .Q(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6498_ (.D(_0131_),
    .CLK(net44),
    .Q(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6499_ (.D(_0132_),
    .CLK(net44),
    .Q(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6500_ (.D(_0133_),
    .CLK(net43),
    .Q(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6501_ (.D(_0134_),
    .CLK(net70),
    .Q(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6502_ (.D(_0135_),
    .CLK(net69),
    .Q(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6503_ (.D(_0136_),
    .CLK(net72),
    .Q(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6504_ (.D(_0137_),
    .CLK(net72),
    .Q(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6505_ (.D(_0138_),
    .CLK(net119),
    .Q(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6506_ (.D(_0139_),
    .CLK(net118),
    .Q(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6507_ (.D(_0140_),
    .CLK(net119),
    .Q(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6508_ (.D(_0141_),
    .CLK(net115),
    .Q(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6509_ (.D(_0142_),
    .CLK(net87),
    .Q(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6510_ (.D(_0143_),
    .CLK(net95),
    .Q(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6511_ (.D(_0144_),
    .CLK(net87),
    .Q(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6512_ (.D(_0145_),
    .CLK(net95),
    .Q(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6513_ (.D(_0146_),
    .CLK(net41),
    .Q(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6514_ (.D(_0147_),
    .CLK(net43),
    .Q(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6515_ (.D(_0148_),
    .CLK(net42),
    .Q(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6516_ (.D(_0149_),
    .CLK(net43),
    .Q(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6517_ (.D(_0150_),
    .CLK(net69),
    .Q(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6518_ (.D(_0151_),
    .CLK(net69),
    .Q(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6519_ (.D(_0152_),
    .CLK(net42),
    .Q(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6520_ (.D(_0153_),
    .CLK(net69),
    .Q(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6521_ (.D(_0154_),
    .CLK(net118),
    .Q(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6522_ (.D(_0155_),
    .CLK(net117),
    .Q(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6523_ (.D(_0156_),
    .CLK(net115),
    .Q(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6524_ (.D(_0157_),
    .CLK(net116),
    .Q(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6525_ (.D(_0158_),
    .CLK(net88),
    .Q(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6526_ (.D(_0159_),
    .CLK(net94),
    .Q(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6527_ (.D(_0160_),
    .CLK(net88),
    .Q(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6528_ (.D(_0161_),
    .CLK(net96),
    .Q(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6529_ (.D(_0162_),
    .CLK(net39),
    .Q(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6530_ (.D(_0163_),
    .CLK(net44),
    .Q(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6531_ (.D(_0164_),
    .CLK(net45),
    .Q(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6532_ (.D(_0165_),
    .CLK(net39),
    .Q(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6533_ (.D(_0166_),
    .CLK(net71),
    .Q(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6534_ (.D(_0167_),
    .CLK(net41),
    .Q(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6535_ (.D(_0168_),
    .CLK(net42),
    .Q(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6536_ (.D(_0169_),
    .CLK(net70),
    .Q(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6537_ (.D(_0170_),
    .CLK(net116),
    .Q(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6538_ (.D(_0171_),
    .CLK(net117),
    .Q(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6539_ (.D(_0172_),
    .CLK(net115),
    .Q(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6540_ (.D(_0173_),
    .CLK(net116),
    .Q(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6541_ (.D(_0174_),
    .CLK(net100),
    .Q(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6542_ (.D(_0175_),
    .CLK(net98),
    .Q(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6543_ (.D(_0176_),
    .CLK(net100),
    .Q(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6544_ (.D(_0177_),
    .CLK(net98),
    .Q(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6545_ (.D(_0178_),
    .CLK(net64),
    .Q(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6546_ (.D(_0179_),
    .CLK(net45),
    .Q(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6547_ (.D(_0180_),
    .CLK(net48),
    .Q(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6548_ (.D(_0181_),
    .CLK(net63),
    .Q(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6549_ (.D(_0182_),
    .CLK(net72),
    .Q(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6550_ (.D(_0183_),
    .CLK(net71),
    .Q(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6551_ (.D(_0184_),
    .CLK(net73),
    .Q(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6552_ (.D(_0185_),
    .CLK(net72),
    .Q(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6553_ (.D(_0186_),
    .CLK(net122),
    .Q(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6554_ (.D(_0187_),
    .CLK(net122),
    .Q(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6555_ (.D(_0188_),
    .CLK(net120),
    .Q(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6556_ (.D(_0189_),
    .CLK(net120),
    .Q(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6557_ (.D(_0190_),
    .CLK(net88),
    .Q(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6558_ (.D(_0191_),
    .CLK(net95),
    .Q(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6559_ (.D(_0192_),
    .CLK(net92),
    .Q(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6560_ (.D(_0193_),
    .CLK(net94),
    .Q(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6561_ (.D(_0194_),
    .CLK(net56),
    .Q(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6562_ (.D(_0195_),
    .CLK(net58),
    .Q(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6563_ (.D(_0196_),
    .CLK(net57),
    .Q(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6564_ (.D(_0197_),
    .CLK(net56),
    .Q(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6565_ (.D(_0198_),
    .CLK(net45),
    .Q(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6566_ (.D(_0199_),
    .CLK(net47),
    .Q(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6567_ (.D(_0200_),
    .CLK(net47),
    .Q(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6568_ (.D(_0201_),
    .CLK(net46),
    .Q(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6569_ (.D(_0202_),
    .CLK(net122),
    .Q(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6570_ (.D(_0203_),
    .CLK(net130),
    .Q(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6571_ (.D(_0204_),
    .CLK(net120),
    .Q(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6572_ (.D(_0205_),
    .CLK(net120),
    .Q(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6573_ (.D(_0206_),
    .CLK(net89),
    .Q(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6574_ (.D(_0207_),
    .CLK(net91),
    .Q(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6575_ (.D(_0208_),
    .CLK(net92),
    .Q(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6576_ (.D(_0209_),
    .CLK(net91),
    .Q(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6577_ (.D(_0210_),
    .CLK(net52),
    .Q(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6578_ (.D(_0211_),
    .CLK(net51),
    .Q(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6579_ (.D(_0212_),
    .CLK(net52),
    .Q(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6580_ (.D(_0213_),
    .CLK(net51),
    .Q(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6581_ (.D(_0214_),
    .CLK(net63),
    .Q(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6582_ (.D(_0215_),
    .CLK(net63),
    .Q(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6583_ (.D(_0216_),
    .CLK(net65),
    .Q(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6584_ (.D(_0217_),
    .CLK(net65),
    .Q(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6585_ (.D(_0218_),
    .CLK(net130),
    .Q(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6586_ (.D(_0219_),
    .CLK(net130),
    .Q(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6587_ (.D(_0220_),
    .CLK(net122),
    .Q(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6588_ (.D(_0221_),
    .CLK(net130),
    .Q(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6589_ (.D(_0222_),
    .CLK(net89),
    .Q(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6590_ (.D(_0223_),
    .CLK(net92),
    .Q(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6591_ (.D(_0224_),
    .CLK(net92),
    .Q(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6592_ (.D(_0225_),
    .CLK(net93),
    .Q(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6593_ (.D(_0226_),
    .CLK(net57),
    .Q(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6594_ (.D(_0227_),
    .CLK(net58),
    .Q(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6595_ (.D(_0228_),
    .CLK(net89),
    .Q(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6596_ (.D(_0229_),
    .CLK(net56),
    .Q(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6597_ (.D(_0230_),
    .CLK(net46),
    .Q(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6598_ (.D(_0231_),
    .CLK(net74),
    .Q(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6599_ (.D(_0232_),
    .CLK(net74),
    .Q(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6600_ (.D(_0233_),
    .CLK(net70),
    .Q(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6601_ (.D(_0234_),
    .CLK(net123),
    .Q(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6602_ (.D(_0235_),
    .CLK(net131),
    .Q(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6603_ (.D(_0236_),
    .CLK(net121),
    .Q(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6604_ (.D(_0237_),
    .CLK(net121),
    .Q(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6605_ (.D(_0238_),
    .CLK(net104),
    .Q(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6606_ (.D(_0239_),
    .CLK(net91),
    .Q(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6607_ (.D(_0240_),
    .CLK(net94),
    .Q(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6608_ (.D(_0241_),
    .CLK(net91),
    .Q(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6609_ (.D(_0242_),
    .CLK(net55),
    .Q(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6610_ (.D(_0243_),
    .CLK(net53),
    .Q(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6611_ (.D(_0244_),
    .CLK(net52),
    .Q(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6612_ (.D(_0245_),
    .CLK(net51),
    .Q(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6613_ (.D(_0246_),
    .CLK(net46),
    .Q(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6614_ (.D(_0247_),
    .CLK(net44),
    .Q(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6615_ (.D(_0248_),
    .CLK(net41),
    .Q(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6616_ (.D(_0249_),
    .CLK(net41),
    .Q(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6617_ (.D(_0250_),
    .CLK(net131),
    .Q(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6618_ (.D(_0251_),
    .CLK(net125),
    .Q(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6619_ (.D(_0252_),
    .CLK(net125),
    .Q(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6620_ (.D(_0253_),
    .CLK(net133),
    .Q(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6621_ (.D(_0254_),
    .CLK(net108),
    .Q(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6622_ (.D(_0255_),
    .CLK(net108),
    .Q(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6623_ (.D(_0256_),
    .CLK(net107),
    .Q(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6624_ (.D(_0257_),
    .CLK(net110),
    .Q(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6625_ (.D(_0258_),
    .CLK(net66),
    .Q(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6626_ (.D(_0259_),
    .CLK(net66),
    .Q(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6627_ (.D(_0260_),
    .CLK(net67),
    .Q(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6628_ (.D(_0261_),
    .CLK(net66),
    .Q(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6629_ (.D(_0262_),
    .CLK(net83),
    .Q(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6630_ (.D(_0263_),
    .CLK(net83),
    .Q(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6631_ (.D(_0264_),
    .CLK(net82),
    .Q(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6632_ (.D(_0265_),
    .CLK(net82),
    .Q(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6633_ (.D(_0266_),
    .CLK(net125),
    .Q(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6634_ (.D(_0267_),
    .CLK(net127),
    .Q(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6635_ (.D(_0268_),
    .CLK(net127),
    .Q(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6636_ (.D(_0269_),
    .CLK(net127),
    .Q(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6637_ (.D(_0270_),
    .CLK(net110),
    .Q(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6638_ (.D(_0271_),
    .CLK(net110),
    .Q(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6639_ (.D(_0272_),
    .CLK(net110),
    .Q(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6640_ (.D(_0273_),
    .CLK(net112),
    .Q(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6641_ (.D(_0274_),
    .CLK(net53),
    .Q(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6642_ (.D(_0275_),
    .CLK(net64),
    .Q(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6643_ (.D(_0276_),
    .CLK(net87),
    .Q(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6644_ (.D(_0277_),
    .CLK(net63),
    .Q(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6645_ (.D(_0278_),
    .CLK(net81),
    .Q(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6646_ (.D(_0279_),
    .CLK(net80),
    .Q(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6647_ (.D(_0280_),
    .CLK(net79),
    .Q(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6648_ (.D(_0281_),
    .CLK(net80),
    .Q(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6649_ (.D(_0282_),
    .CLK(net123),
    .Q(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6650_ (.D(_0283_),
    .CLK(net123),
    .Q(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6651_ (.D(_0284_),
    .CLK(net121),
    .Q(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6652_ (.D(_0285_),
    .CLK(net121),
    .Q(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6653_ (.D(_0286_),
    .CLK(net107),
    .Q(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6654_ (.D(_0287_),
    .CLK(net107),
    .Q(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6655_ (.D(_0288_),
    .CLK(net105),
    .Q(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6656_ (.D(_0289_),
    .CLK(net107),
    .Q(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6657_ (.D(_0290_),
    .CLK(net54),
    .Q(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6658_ (.D(_0291_),
    .CLK(net59),
    .Q(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6659_ (.D(_0292_),
    .CLK(net60),
    .Q(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6660_ (.D(_0293_),
    .CLK(net54),
    .Q(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6661_ (.D(_0294_),
    .CLK(net81),
    .Q(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6662_ (.D(_0295_),
    .CLK(net80),
    .Q(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6663_ (.D(_0296_),
    .CLK(net79),
    .Q(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6664_ (.D(_0297_),
    .CLK(net79),
    .Q(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6665_ (.D(_0298_),
    .CLK(net132),
    .Q(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6666_ (.D(_0299_),
    .CLK(net133),
    .Q(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6667_ (.D(_0300_),
    .CLK(net131),
    .Q(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6668_ (.D(_0301_),
    .CLK(net135),
    .Q(\mod.registers.r12[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6669_ (.D(_0302_),
    .CLK(net105),
    .Q(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6670_ (.D(_0303_),
    .CLK(net111),
    .Q(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6671_ (.D(_0304_),
    .CLK(net111),
    .Q(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6672_ (.D(_0305_),
    .CLK(net111),
    .Q(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6673_ (.D(_0306_),
    .CLK(net59),
    .Q(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6674_ (.D(_0307_),
    .CLK(net60),
    .Q(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6675_ (.D(_0308_),
    .CLK(net87),
    .Q(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6676_ (.D(_0309_),
    .CLK(net59),
    .Q(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6677_ (.D(_0310_),
    .CLK(net83),
    .Q(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6678_ (.D(_0311_),
    .CLK(net83),
    .Q(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6679_ (.D(_0312_),
    .CLK(net82),
    .Q(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6680_ (.D(_0313_),
    .CLK(net82),
    .Q(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6681_ (.D(_0314_),
    .CLK(net133),
    .Q(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6682_ (.D(_0315_),
    .CLK(net133),
    .Q(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6683_ (.D(_0316_),
    .CLK(net126),
    .Q(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6684_ (.D(_0317_),
    .CLK(net134),
    .Q(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6685_ (.D(_0318_),
    .CLK(net102),
    .Q(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6686_ (.D(_0319_),
    .CLK(net98),
    .Q(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6687_ (.D(_0320_),
    .CLK(net94),
    .Q(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6688_ (.D(_0321_),
    .CLK(net105),
    .Q(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6689_ (.D(_0322_),
    .CLK(net54),
    .Q(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6690_ (.D(_0323_),
    .CLK(net40),
    .Q(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6691_ (.D(_0324_),
    .CLK(net39),
    .Q(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6692_ (.D(_0325_),
    .CLK(net53),
    .Q(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6693_ (.D(_0326_),
    .CLK(net76),
    .Q(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6694_ (.D(_0327_),
    .CLK(net74),
    .Q(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6695_ (.D(_0328_),
    .CLK(net76),
    .Q(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6696_ (.D(_0329_),
    .CLK(net76),
    .Q(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6697_ (.D(_0330_),
    .CLK(net126),
    .Q(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6698_ (.D(_0331_),
    .CLK(net126),
    .Q(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6699_ (.D(_0332_),
    .CLK(net125),
    .Q(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6700_ (.D(_0333_),
    .CLK(net127),
    .Q(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6701_ (.D(_0334_),
    .CLK(net106),
    .Q(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6702_ (.D(_0335_),
    .CLK(net105),
    .Q(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6703_ (.D(_0336_),
    .CLK(net103),
    .Q(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6704_ (.D(_0337_),
    .CLK(net106),
    .Q(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6705_ (.D(_0338_),
    .CLK(net53),
    .Q(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6706_ (.D(_0339_),
    .CLK(net39),
    .Q(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6707_ (.D(_0340_),
    .CLK(net40),
    .Q(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6708_ (.D(_0341_),
    .CLK(net51),
    .Q(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6709_ (.D(_0342_),
    .CLK(net77),
    .Q(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6710_ (.D(_0343_),
    .CLK(net75),
    .Q(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6711_ (.D(_0344_),
    .CLK(net76),
    .Q(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6712_ (.D(_0345_),
    .CLK(net74),
    .Q(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6713_ (.D(_0000_),
    .SETN(_0004_),
    .CLK(net201),
    .Q(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6714_ (.D(_0001_),
    .SETN(_0005_),
    .CLK(net201),
    .Q(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _6715_ (.D(_0002_),
    .SETN(_0006_),
    .CLK(net201),
    .Q(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6716_ (.D(_0346_),
    .CLK(net189),
    .Q(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6717_ (.D(_0347_),
    .CLK(net184),
    .Q(\mod.valid1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6718_ (.D(_0348_),
    .CLK(net148),
    .Q(\mod.pc0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6719_ (.D(_0349_),
    .CLK(net147),
    .Q(\mod.pc0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6720_ (.D(_0350_),
    .CLK(net142),
    .Q(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6721_ (.D(_0351_),
    .CLK(net143),
    .Q(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6722_ (.D(_0352_),
    .CLK(net144),
    .Q(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6723_ (.D(_0353_),
    .CLK(net148),
    .Q(\mod.pc0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6724_ (.D(_0354_),
    .CLK(net144),
    .Q(\mod.pc0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6725_ (.D(_0355_),
    .CLK(net142),
    .Q(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6726_ (.D(_0356_),
    .CLK(net150),
    .Q(\mod.pc0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6727_ (.D(_0357_),
    .CLK(net144),
    .Q(\mod.pc0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6728_ (.D(_0358_),
    .CLK(net148),
    .Q(\mod.pc0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6729_ (.D(_0359_),
    .CLK(net141),
    .Q(\mod.pc0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6730_ (.D(_0360_),
    .CLK(net141),
    .Q(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6731_ (.D(_0361_),
    .CLK(net141),
    .Q(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6732_ (.D(_0362_),
    .CLK(net152),
    .Q(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6733_ (.D(_0363_),
    .CLK(net149),
    .Q(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6734_ (.D(_0364_),
    .CLK(net153),
    .Q(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6735_ (.D(_0365_),
    .CLK(net152),
    .Q(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6736_ (.D(_0366_),
    .CLK(net153),
    .Q(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6737_ (.D(_0367_),
    .CLK(net151),
    .Q(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6738_ (.D(_0368_),
    .CLK(net151),
    .Q(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6739_ (.D(_0369_),
    .CLK(net151),
    .Q(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6740_ (.D(_0370_),
    .CLK(net149),
    .Q(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6741_ (.D(_0371_),
    .CLK(net149),
    .Q(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6742_ (.D(_0372_),
    .CLK(net149),
    .Q(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6743_ (.D(_0373_),
    .CLK(net144),
    .Q(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6744_ (.D(_0374_),
    .CLK(net150),
    .Q(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6745_ (.D(_0375_),
    .CLK(net145),
    .Q(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6746_ (.D(_0376_),
    .CLK(net186),
    .Q(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6747_ (.D(_0377_),
    .CLK(net187),
    .Q(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6748_ (.D(_0378_),
    .CLK(net187),
    .Q(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6749_ (.D(_0379_),
    .CLK(net188),
    .Q(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6750_ (.D(_0380_),
    .CLK(net187),
    .Q(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6751_ (.D(_0381_),
    .CLK(net186),
    .Q(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6752_ (.D(_0382_),
    .CLK(net186),
    .Q(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6753_ (.D(_0383_),
    .CLK(net151),
    .Q(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6754_ (.D(_0384_),
    .CLK(net186),
    .Q(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6755_ (.D(_0385_),
    .CLK(net153),
    .Q(\mod.pc_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6756_ (.D(_0386_),
    .CLK(net187),
    .Q(\mod.pc_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6757_ (.D(_0387_),
    .CLK(net152),
    .Q(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6758_ (.D(_0388_),
    .CLK(net155),
    .Q(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6759_ (.D(_0389_),
    .CLK(net180),
    .Q(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6760_ (.D(_0390_),
    .CLK(net175),
    .Q(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6761_ (.D(_0391_),
    .CLK(net175),
    .Q(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6762_ (.D(_0392_),
    .CLK(net176),
    .Q(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6763_ (.D(_0393_),
    .CLK(net175),
    .Q(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6764_ (.D(_0394_),
    .CLK(net170),
    .Q(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6765_ (.D(_0395_),
    .CLK(net173),
    .Q(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6766_ (.D(_0396_),
    .CLK(net173),
    .Q(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6767_ (.D(_0397_),
    .CLK(net173),
    .Q(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6768_ (.D(_0398_),
    .CLK(net174),
    .Q(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6769_ (.D(_0399_),
    .CLK(net174),
    .Q(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6770_ (.D(_0400_),
    .CLK(net173),
    .Q(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6771_ (.D(_0401_),
    .CLK(net168),
    .Q(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6772_ (.D(_0402_),
    .CLK(net168),
    .Q(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6773_ (.D(_0403_),
    .CLK(net167),
    .Q(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6774_ (.D(_0404_),
    .CLK(net167),
    .Q(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6775_ (.D(_0405_),
    .CLK(net167),
    .Q(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6776_ (.D(_0406_),
    .CLK(net165),
    .Q(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6777_ (.D(_0407_),
    .CLK(net168),
    .Q(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6778_ (.D(_0408_),
    .CLK(net166),
    .Q(\mod.instr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6779_ (.D(_0409_),
    .CLK(net166),
    .Q(\mod.instr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6780_ (.D(_0007_),
    .CLK(net167),
    .Q(\mod.instr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6781_ (.D(_0008_),
    .CLK(net182),
    .Q(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6782_ (.D(_0009_),
    .CLK(net161),
    .Q(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6783_ (.D(_0010_),
    .CLK(net160),
    .Q(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6784_ (.D(_0011_),
    .CLK(net160),
    .Q(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6785_ (.D(_0012_),
    .CLK(net175),
    .Q(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6786_ (.D(_0013_),
    .CLK(net170),
    .Q(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6787_ (.D(_0014_),
    .CLK(net172),
    .Q(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6788_ (.D(_0015_),
    .CLK(net172),
    .Q(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6789_ (.D(_0016_),
    .CLK(net160),
    .Q(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6790_ (.D(_0017_),
    .CLK(net158),
    .Q(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6791_ (.D(_0018_),
    .CLK(net159),
    .Q(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6792_ (.D(_0019_),
    .CLK(net158),
    .Q(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6793_ (.D(_0020_),
    .CLK(net158),
    .Q(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6794_ (.D(_0021_),
    .CLK(net158),
    .Q(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6795_ (.D(_0022_),
    .CLK(net165),
    .Q(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6796_ (.D(_0023_),
    .CLK(net166),
    .Q(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6797_ (.D(_0024_),
    .CLK(net165),
    .Q(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6798_ (.D(_0025_),
    .CLK(net165),
    .Q(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6799_ (.D(_0026_),
    .CLK(net132),
    .Q(\mod.instr_2[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6800_ (.D(_0027_),
    .CLK(net169),
    .Q(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6801_ (.D(_0028_),
    .CLK(net171),
    .Q(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6802_ (.D(_0029_),
    .CLK(net170),
    .Q(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6803_ (.D(_0030_),
    .CLK(net180),
    .Q(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6804_ (.D(_0031_),
    .CLK(net181),
    .Q(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6805_ (.D(_0032_),
    .CLK(net181),
    .Q(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6806_ (.D(_0033_),
    .CLK(net162),
    .Q(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6807_ (.D(_0034_),
    .CLK(net162),
    .Q(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6808_ (.D(_0035_),
    .CLK(net162),
    .Q(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6809_ (.D(_0036_),
    .CLK(net162),
    .Q(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6810_ (.D(_0037_),
    .CLK(net157),
    .Q(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6811_ (.D(_0038_),
    .CLK(net157),
    .Q(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6812_ (.D(_0039_),
    .CLK(net157),
    .Q(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6813_ (.D(_0040_),
    .CLK(net157),
    .Q(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6814_ (.D(_0041_),
    .CLK(net147),
    .Q(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6815_ (.D(_0042_),
    .CLK(net147),
    .Q(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6816_ (.D(_0043_),
    .CLK(net147),
    .Q(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0044_),
    .CLK(net161),
    .Q(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0045_),
    .CLK(net160),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0046_),
    .CLK(net180),
    .Q(\mod.ri_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0047_),
    .CLK(net182),
    .Q(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0048_),
    .CLK(net180),
    .Q(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0049_),
    .CLK(net182),
    .Q(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0050_),
    .CLK(net184),
    .Q(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0051_),
    .CLK(net182),
    .Q(\mod.rd_3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0052_),
    .CLK(net193),
    .Q(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0053_),
    .CLK(net193),
    .Q(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0054_),
    .CLK(net191),
    .Q(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0055_),
    .CLK(net191),
    .Q(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6829_ (.D(_0056_),
    .CLK(net191),
    .Q(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6830_ (.D(_0057_),
    .CLK(net192),
    .Q(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6831_ (.D(_0058_),
    .CLK(net192),
    .Q(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6832_ (.D(_0059_),
    .CLK(net192),
    .Q(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6833_ (.D(_0060_),
    .CLK(net171),
    .Q(\mod.ldr_hzd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6834_ (.D(_0061_),
    .CLK(net170),
    .Q(\mod.ldr_hzd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6835_ (.D(_0062_),
    .CLK(net171),
    .Q(\mod.ldr_hzd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6836_ (.D(_0063_),
    .CLK(net172),
    .Q(\mod.ldr_hzd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6837_ (.D(_0064_),
    .CLK(net183),
    .Q(\mod.ldr_hzd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6838_ (.D(_0065_),
    .CLK(net183),
    .Q(\mod.ldr_hzd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6839_ (.D(_0066_),
    .CLK(net191),
    .Q(\mod.ldr_hzd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6840_ (.D(_0067_),
    .CLK(net183),
    .Q(\mod.ldr_hzd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6841_ (.D(_0068_),
    .CLK(net212),
    .Q(\mod.des.des_dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6842_ (.D(_0069_),
    .CLK(net212),
    .Q(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6843_ (.D(_0070_),
    .CLK(net211),
    .Q(\mod.des.des_dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6844_ (.D(_0071_),
    .CLK(net211),
    .Q(\mod.des.des_dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6845_ (.D(_0072_),
    .CLK(net207),
    .Q(\mod.des.des_dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6846_ (.D(_0073_),
    .CLK(net205),
    .Q(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6847_ (.D(_0074_),
    .CLK(net205),
    .Q(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6848_ (.D(_0075_),
    .CLK(net205),
    .Q(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6849_ (.D(_0076_),
    .CLK(net208),
    .Q(\mod.des.des_dout[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6850_ (.D(_0077_),
    .CLK(net209),
    .Q(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6851_ (.D(_0078_),
    .CLK(net211),
    .Q(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6852_ (.D(_0079_),
    .CLK(net209),
    .Q(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6853_ (.D(_0080_),
    .CLK(net211),
    .Q(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6854_ (.D(_0081_),
    .CLK(net135),
    .Q(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6855_ (.D(_0082_),
    .CLK(net134),
    .Q(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6856_ (.D(_0083_),
    .CLK(net134),
    .Q(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6857_ (.D(_0084_),
    .CLK(net135),
    .Q(\mod.registers.r15[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6858_ (.D(_0085_),
    .CLK(net102),
    .Q(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6859_ (.D(_0086_),
    .CLK(net102),
    .Q(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6860_ (.D(_0087_),
    .CLK(net103),
    .Q(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6861_ (.D(_0088_),
    .CLK(net102),
    .Q(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6862_ (.D(_0089_),
    .CLK(net59),
    .Q(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6863_ (.D(_0090_),
    .CLK(net57),
    .Q(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6864_ (.D(_0091_),
    .CLK(net89),
    .Q(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6865_ (.D(_0092_),
    .CLK(net56),
    .Q(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6866_ (.D(_0093_),
    .CLK(net75),
    .Q(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6867_ (.D(_0094_),
    .CLK(net75),
    .Q(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6868_ (.D(_0095_),
    .CLK(net46),
    .Q(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6869_ (.D(_0096_),
    .CLK(net79),
    .Q(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6870_ (.D(_0097_),
    .CLK(net209),
    .Q(\mod.des.des_dout[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6871_ (.D(_0098_),
    .CLK(net208),
    .Q(\mod.des.des_dout[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6872_ (.D(_0099_),
    .CLK(net208),
    .Q(\mod.des.des_dout[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6873_ (.D(_0100_),
    .CLK(net208),
    .Q(\mod.des.des_dout[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6874_ (.D(_0101_),
    .CLK(net205),
    .Q(\mod.des.des_dout[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6875_ (.D(_0102_),
    .CLK(net206),
    .Q(\mod.des.des_dout[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6876_ (.D(_0103_),
    .CLK(net206),
    .Q(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6877_ (.D(_0104_),
    .CLK(net206),
    .Q(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6878_ (.D(_0105_),
    .CLK(net198),
    .Q(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6879_ (.D(_0106_),
    .CLK(net202),
    .Q(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6880_ (.D(_0107_),
    .CLK(net202),
    .Q(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6881_ (.D(_0108_),
    .CLK(net202),
    .Q(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6882_ (.D(_0109_),
    .CLK(net212),
    .Q(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6883_ (.D(_0110_),
    .CLK(net204),
    .Q(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6884_ (.D(_0111_),
    .CLK(net202),
    .Q(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6885_ (.D(_0112_),
    .CLK(net204),
    .Q(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6886_ (.D(_0113_),
    .CLK(net204),
    .Q(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6887_ (.D(_0114_),
    .CLK(net198),
    .Q(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6888_ (.D(_0115_),
    .CLK(net198),
    .Q(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6889_ (.D(_0116_),
    .CLK(net199),
    .Q(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6890_ (.D(_0117_),
    .CLK(net198),
    .Q(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6891_ (.D(_0118_),
    .CLK(net200),
    .Q(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6892_ (.D(_0119_),
    .CLK(net203),
    .Q(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6893_ (.D(_0120_),
    .CLK(net200),
    .Q(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_295 (.ZN(net295));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_296 (.ZN(net296));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_297 (.ZN(net297));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_331 (.ZN(net331));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_332 (.ZN(net332));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_333 (.ZN(net333));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_334 (.ZN(net334));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_335 (.ZN(net335));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_336 (.ZN(net336));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_337 (.ZN(net337));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_338 (.ZN(net338));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_339 (.ZN(net339));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_340 (.ZN(net340));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_341 (.ZN(net341));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_342 (.ZN(net342));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_343 (.ZN(net343));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_344 (.ZN(net344));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_345 (.ZN(net345));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_346 (.ZN(net346));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_347 (.ZN(net347));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_348 (.ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_349 (.ZN(net349));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_350 (.ZN(net350));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_351 (.ZN(net351));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_352 (.ZN(net352));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_353 (.ZN(net353));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_354 (.ZN(net354));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_355 (.ZN(net355));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_356 (.ZN(net356));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_357 (.ZN(net357));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_358 (.ZN(net358));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_359 (.ZN(net359));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_360 (.ZN(net360));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_361 (.ZN(net361));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_362 (.ZN(net362));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_363 (.ZN(net363));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_364 (.ZN(net364));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_365 (.ZN(net365));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_366 (.ZN(net366));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_367 (.ZN(net367));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_368 (.ZN(net368));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_369 (.ZN(net369));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_370 (.ZN(net370));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_371 (.ZN(net371));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_372 (.ZN(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(io_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input11 (.I(io_in[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input12 (.I(io_in[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(io_in[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_in[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(io_in[5]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(io_in[6]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(io_in[7]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(io_in[8]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(io_in[9]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout40 (.I(net50),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout42 (.I(net49),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net49),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net48),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net68),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net55),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net55),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net62),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net61),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net61),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net67),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net86),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net73),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net73),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net78),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout74 (.I(net77),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net77),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net85),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net84),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net84),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout82 (.I(net84),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net140),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout87 (.I(net90),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net90),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout89 (.I(net97),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout90 (.I(net97),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net93),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout92 (.I(net96),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net96),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout95 (.I(net96),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net97),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout97 (.I(net101),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net101),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net101),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout101 (.I(net114),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout102 (.I(net104),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net113),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net109),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net109),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout107 (.I(net109),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net112),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net111),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout114 (.I(net139),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout115 (.I(net119),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout117 (.I(net118),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout119 (.I(net138),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout120 (.I(net124),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout121 (.I(net124),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout122 (.I(net124),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net129),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout125 (.I(net128),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net128),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout127 (.I(net129),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net137),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout130 (.I(net132),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net136),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout133 (.I(net134),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout134 (.I(net135),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout135 (.I(net136),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net138),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout138 (.I(net139),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net197),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout141 (.I(net143),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout143 (.I(net146),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net146),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net156),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net155),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net154),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout151 (.I(net154),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout152 (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout153 (.I(net154),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout154 (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout155 (.I(net156),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net196),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout157 (.I(net196),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout158 (.I(net159),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout159 (.I(net164),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout160 (.I(net163),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout161 (.I(net163),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout162 (.I(net164),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout163 (.I(net164),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout164 (.I(net179),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout165 (.I(net166),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout166 (.I(net169),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout167 (.I(net169),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout168 (.I(net169),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net178),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net171),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout171 (.I(net172),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout172 (.I(net177),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout173 (.I(net176),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout174 (.I(net176),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout176 (.I(net177),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout177 (.I(net178),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout178 (.I(net179),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout179 (.I(net195),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout180 (.I(net181),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout181 (.I(net185),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout182 (.I(net183),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout183 (.I(net185),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout184 (.I(net185),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout185 (.I(net190),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout186 (.I(net188),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout187 (.I(net189),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout188 (.I(net189),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout189 (.I(net190),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout190 (.I(net194),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout191 (.I(net193),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout192 (.I(net193),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout193 (.I(net194),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout194 (.I(net195),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout195 (.I(net196),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout196 (.I(net197),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout197 (.I(\mod.clk ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout198 (.I(net199),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net200),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout200 (.I(net215),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout201 (.I(net215),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout202 (.I(net203),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout203 (.I(net204),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout204 (.I(net214),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout205 (.I(net206),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout206 (.I(net207),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout207 (.I(net210),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout208 (.I(net210),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout209 (.I(net210),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout210 (.I(net213),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout211 (.I(net212),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout212 (.I(net213),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout213 (.I(net214),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net215),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net1),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__RN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__D (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__D (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__D (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__D (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__C (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__C1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__C1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__B1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__B1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__B1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__C1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__C1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__B1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__B1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__B1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__B1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__B1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__C1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A3 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__B (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__C (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__I0 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__B (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__I1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__S (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__S (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__I (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__B (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__B (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__B1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__B1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__B1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__A4 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__B2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__I (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__C1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__I (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__B1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__B1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__B1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__I (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__C2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__C2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__B1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__B1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__B1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__B1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__B1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__I (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__B1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__B1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__C1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__B1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__C1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__B1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A3 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__B (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__B (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__B (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__B (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__I1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__I0 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__B1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__B1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__B1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__B1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__B1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__B2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__B (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__I0 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__I1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__B1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__B1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__C1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__B1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__B1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A3 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__B1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__B1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__B1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__B1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__C1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__B1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__C1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__B1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__B1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__B1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__B1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A3 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__B (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A3 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__B (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I0 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__B (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__I (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__B (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__B (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A3 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A3 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A3 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__B2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__C (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A4 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A3 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A3 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__S (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A3 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A3 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__B1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__C2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__C2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__C (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__B2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A3 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__B (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A3 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__B2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__C (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A3 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__C (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__I0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__B1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__B2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A3 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__B (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__B1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__B2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I0 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A3 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__B (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A4 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A4 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A3 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A3 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__I (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__I (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__I1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__C (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A4 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A4 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__B2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A3 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I3 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__B (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__B (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A3 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__B2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A3 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__B (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A3 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A3 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__I (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A3 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A3 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__B2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A3 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__B1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__B2 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A3 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__B (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__B (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__B2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__C (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__B1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__B1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__B1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__B1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__B1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__B1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__B1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__B1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__B1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__B1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__B1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__B1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__B (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__B1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__B1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__B1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__B1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__C2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__C2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__C2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__C2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__C1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__C1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__B1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__B1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__B1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__B1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__B1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A3 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__B (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__B (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__B (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A3 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__B (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__B2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I3 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__C (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A3 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__B1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__B1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__C1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__C1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__C1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__C1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A3 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__B1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__B1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A3 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A3 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A3 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I0 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I0 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__B (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__C1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__B1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A3 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A3 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A3 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A3 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__B (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A3 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__B1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__B (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I3 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__B (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I0 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__C1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__B1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__B1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__B1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__B1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__B1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__B1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__B1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__B1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__C1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__B1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__B2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__B1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__C1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__B1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__B1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__C1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__B1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__B1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__I (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A3 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__B (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__I (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__I (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__B (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__B1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__B2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A3 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I3 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I3 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__I (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__I (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A3 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A3 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A3 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__B (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I0 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A3 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I0 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__I (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__B (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__I (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__B (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__I (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__B (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__I (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__I (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__I (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__B1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__B2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A3 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A3 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__B (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I0 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A3 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I0 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I0 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A3 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__B (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__B (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__B2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__B (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__C (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__S1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__I (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__B2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A3 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__B2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__C (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__S1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__S1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__S (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__S0 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__S0 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__S (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__S1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A3 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__C (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__B (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A3 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A3 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__B1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A3 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__I (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__I (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__I (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__B1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__B (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__B (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__B (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__C (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__S (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__C (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__S1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__B2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__S (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__I (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__B (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__C (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I3 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__B (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I0 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__S0 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__S1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__S0 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__B (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__S (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__S (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__S (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I0 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__I0 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__I1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__B (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I0 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__S (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__B2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__B (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__C (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__B1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__B (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__I (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__I (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__B (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__B (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__B2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__B2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__B (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__B (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__B (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__B (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__B (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__B1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__I (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__B1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__C (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__C (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__C (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__C (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__C (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__S (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__S (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__S0 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__S0 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__S0 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__S (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__C (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__C (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__S1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__B (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__B2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A4 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A3 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A3 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__S (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__S0 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__B (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__C (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__S (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__S (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A3 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__B2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__C (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__C (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__I (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__B2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__C (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__B (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__I (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__C (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__B (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__B (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__B (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__I (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__C (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__B (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__C (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A3 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__B (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__C (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__C (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A3 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I0 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I3 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I0 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__C (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__B (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__B (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A3 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I0 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I0 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I3 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__B1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__B1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__B2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__B2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__B (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__B (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__B (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I0 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__B1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__B1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__B2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__C (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__B2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A3 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I0 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__B1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I0 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I0 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__C (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__C (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__C (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A3 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__I1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__B1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A3 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__C (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__B1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__C (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__B1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__B2 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__C (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A4 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__B1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A4 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A3 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__B (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__C (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A4 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A3 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A3 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__B1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__B (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__B (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__C (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__C (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__B (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__C (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A3 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__B (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__B (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__C (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__B (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__B1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A4 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I0 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A3 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__C2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I3 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__S0 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__S0 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__S1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__S1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A4 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I0 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A3 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__C2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I3 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A3 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__B2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__B2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A3 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__C2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__B2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A4 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__B2 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__C1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__B (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__B1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__B1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__C1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__C1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__C1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__C1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A4 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__B2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__C1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__B1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__B1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__B1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__B1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__B1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__C (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__B2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__B1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A3 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__C (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__B2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__S (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__C (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__I (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__B1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__B1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__B1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__B2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__B (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__B (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__B (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__B2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__B (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__B (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__C (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__I (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__B (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A3 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__C (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__B1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__I (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__B1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__B2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__B1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__B2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__B2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__B2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__C (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__B1 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A3 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A2 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__C (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__B1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__B (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__B2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__C (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A3 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__B1 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__B2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__C (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__S (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__B2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__B (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__B (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A3 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A3 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__B1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B1 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I1 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A3 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__B1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__I (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A3 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__B (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__I (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__B (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__B (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__B (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__B (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__B (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__B (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__B (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__B1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__B1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__B1 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__I (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__I (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__B1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__B1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__I (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__I (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A2 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__I (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__I (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__I (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__I (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__I (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__I (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__I (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__I (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__I (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__I (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__I (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__I (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__I (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__I (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__I (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__I (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__I (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__I (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A3 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__I (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__I (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A3 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__I (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A3 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__I (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__I (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__I (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A3 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__B (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__B (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__B (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__I (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__B (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__B (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__B (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__B (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__C (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__C (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A2 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__B (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__B (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__B (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__C (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__C (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__C (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__C (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__C (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A4 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__I (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__I (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__I (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__I (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__I (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__B (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__I (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__I (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__I (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__I (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__B2 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__I (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__I (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__I (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__B2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__B2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__B2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__B2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B1 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__C (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__C (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__C (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__C (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__C (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__I (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__B1 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__B1 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__B1 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B1 (.I(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__B (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__B (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__B (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__B (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__B (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__B (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A4 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A2 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A3 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__B (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__B (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__B (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__I (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__I (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__B2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__B2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__S (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__S (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__S (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__S (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__S (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__I (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__I (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__I (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__I (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__I (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__I (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__S (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__I (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__I (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__S (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__S (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__S (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__S (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__S (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__S (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__S (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__S (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__I (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__I (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__S (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__S (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__S (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__I (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__S (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__S (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__S (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__S (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__S (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__S (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__S (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__S (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__B (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__I (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__I (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__B (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__I (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A2 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__C (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__I (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A1 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__B (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A3 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__B (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A2 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A2 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__B (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__B (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__I (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__B1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__I (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__I (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__C (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__I (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__I (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__I (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__I (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__I (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__B1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__B1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__B1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__B (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__I (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__I (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A3 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__B (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__B (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__B (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__B1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__I (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__B1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__B1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__I (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__I (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__B1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__B1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__B1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A3 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__B1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__B1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__B1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__B2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I2 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__I0 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__B (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__I (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__I (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__I (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A2 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__I (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A3 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A3 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__B1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__I (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A3 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__B1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__I (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B1 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__B1 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__C1 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__I (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A2 (.I(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__I (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__B1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__I (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__I (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__B1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A3 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A3 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__B1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__B1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__B1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__B1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__B1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__C2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__I (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__C1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__I (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__I (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A3 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__I (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__B1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__A1 (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__I (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__I (.I(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__A2 (.I(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__I (.I(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A3 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A1 (.I(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__I0 (.I(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__I0 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I0 (.I(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__I0 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I0 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I0 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I0 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__I0 (.I(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I0 (.I(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__I0 (.I(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__I0 (.I(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__I1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__I (.I(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I0 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__I (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__I (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B2 (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__B2 (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__I (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B2 (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__B2 (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__I (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__B2 (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__I (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__B2 (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__I (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__B2 (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__I (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__B2 (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__I (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__B2 (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__I (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__B2 (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I (.I(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__B2 (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__B2 (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__I (.I(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__B2 (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I (.I(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__C (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__B (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__I (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A1 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__I (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__I0 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__B2 (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__I (.I(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__B (.I(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I0 (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I1 (.I(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__I (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__I (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__I (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__B (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__B (.I(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__I (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__I (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__I (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__I (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__I (.I(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__I (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__I (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__B2 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__B2 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__B2 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__B2 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A1 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__B2 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B2 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__B2 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__B2 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B2 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__B2 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__B2 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A1 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__B2 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__B2 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__B2 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__B2 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__B2 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B2 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__B2 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__C2 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__B2 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B2 (.I(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B2 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__B2 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__B2 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__B2 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__B2 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__C2 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__C2 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A1 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__B2 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__C2 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__B2 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__B2 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__B2 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__B2 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__C2 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__B2 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B2 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__B2 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__B2 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B2 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B2 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__B2 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__B2 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B2 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__B2 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__B2 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B2 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__B2 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B2 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__B2 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__B2 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__B2 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__C2 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B2 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A3 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B2 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__C1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__B2 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__C1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B2 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__B2 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__C1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__C1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__C2 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__B2 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__C1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A3 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__B2 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__B2 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B2 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__C2 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__B2 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__C1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__B2 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B2 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__B2 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__B2 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__B2 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__B2 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B2 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B2 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__B2 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__B2 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__B2 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B2 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__B2 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B2 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A3 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B2 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__B2 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__B2 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__B2 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B2 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__B2 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A1 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B2 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B2 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__B2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__B2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__B2 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__B2 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__B2 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A3 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B2 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__B2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__B2 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__B2 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__B2 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__B2 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__B2 (.I(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__B2 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__B2 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__C2 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__C2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__B2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__B2 (.I(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B2 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__B2 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B2 (.I(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__B2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__B2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__B2 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__B2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__B2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__B2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__B2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__B2 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__B2 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__B2 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B2 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__B2 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__C2 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A3 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B2 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B2 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__B2 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B2 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__B2 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B2 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__B2 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__B2 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B2 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__C2 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__B2 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__B2 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__B2 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__C2 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__B2 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B2 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__B2 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__B2 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__B2 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__B2 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B2 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B2 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__C2 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B2 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__C2 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__C2 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__B2 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B2 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__B2 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__B2 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__B2 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__B2 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__B2 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__C2 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__B2 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__B2 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__B2 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B2 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B2 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__C2 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B2 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__B2 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__B2 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B2 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__C2 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__C2 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__B2 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B2 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__B2 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__B2 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__B2 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__B2 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__B2 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__B2 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__B2 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__B2 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__I (.I(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__CLK (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__A1 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__CLK (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__CLK (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__CLK (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__CLK (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__CLK (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__CLK (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__CLK (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__CLK (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout166_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__CLK (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__CLK (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__CLK (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__CLK (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout173_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout174_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout169_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout178_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout182_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout179_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout199_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__CLK (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__CLK (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__CLK (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout205_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout206_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1043 ();
 assign io_oeb[0] = net216;
 assign io_oeb[10] = net226;
 assign io_oeb[11] = net227;
 assign io_oeb[12] = net228;
 assign io_oeb[13] = net229;
 assign io_oeb[14] = net230;
 assign io_oeb[15] = net231;
 assign io_oeb[16] = net232;
 assign io_oeb[17] = net233;
 assign io_oeb[18] = net234;
 assign io_oeb[19] = net235;
 assign io_oeb[1] = net217;
 assign io_oeb[20] = net236;
 assign io_oeb[21] = net237;
 assign io_oeb[22] = net238;
 assign io_oeb[23] = net239;
 assign io_oeb[24] = net240;
 assign io_oeb[25] = net241;
 assign io_oeb[26] = net242;
 assign io_oeb[27] = net243;
 assign io_oeb[28] = net244;
 assign io_oeb[29] = net245;
 assign io_oeb[2] = net218;
 assign io_oeb[30] = net246;
 assign io_oeb[31] = net247;
 assign io_oeb[32] = net248;
 assign io_oeb[33] = net249;
 assign io_oeb[34] = net250;
 assign io_oeb[35] = net251;
 assign io_oeb[36] = net252;
 assign io_oeb[37] = net253;
 assign io_oeb[3] = net219;
 assign io_oeb[4] = net220;
 assign io_oeb[5] = net221;
 assign io_oeb[6] = net222;
 assign io_oeb[7] = net223;
 assign io_oeb[8] = net224;
 assign io_oeb[9] = net225;
 assign io_out[0] = net254;
 assign io_out[10] = net264;
 assign io_out[11] = net265;
 assign io_out[12] = net266;
 assign io_out[13] = net267;
 assign io_out[14] = net268;
 assign io_out[15] = net269;
 assign io_out[16] = net270;
 assign io_out[17] = net271;
 assign io_out[18] = net272;
 assign io_out[1] = net255;
 assign io_out[2] = net256;
 assign io_out[3] = net257;
 assign io_out[4] = net258;
 assign io_out[5] = net259;
 assign io_out[6] = net260;
 assign io_out[7] = net261;
 assign io_out[8] = net262;
 assign io_out[9] = net263;
 assign la_data_out[0] = net273;
 assign la_data_out[10] = net283;
 assign la_data_out[11] = net284;
 assign la_data_out[12] = net285;
 assign la_data_out[13] = net286;
 assign la_data_out[14] = net287;
 assign la_data_out[15] = net288;
 assign la_data_out[16] = net289;
 assign la_data_out[17] = net290;
 assign la_data_out[18] = net291;
 assign la_data_out[19] = net292;
 assign la_data_out[1] = net274;
 assign la_data_out[20] = net293;
 assign la_data_out[21] = net294;
 assign la_data_out[22] = net295;
 assign la_data_out[23] = net296;
 assign la_data_out[24] = net297;
 assign la_data_out[25] = net298;
 assign la_data_out[26] = net299;
 assign la_data_out[27] = net300;
 assign la_data_out[28] = net301;
 assign la_data_out[29] = net302;
 assign la_data_out[2] = net275;
 assign la_data_out[30] = net303;
 assign la_data_out[31] = net304;
 assign la_data_out[32] = net305;
 assign la_data_out[33] = net306;
 assign la_data_out[34] = net307;
 assign la_data_out[35] = net308;
 assign la_data_out[36] = net309;
 assign la_data_out[37] = net310;
 assign la_data_out[38] = net311;
 assign la_data_out[39] = net312;
 assign la_data_out[3] = net276;
 assign la_data_out[40] = net313;
 assign la_data_out[41] = net314;
 assign la_data_out[42] = net315;
 assign la_data_out[43] = net316;
 assign la_data_out[44] = net317;
 assign la_data_out[45] = net318;
 assign la_data_out[46] = net319;
 assign la_data_out[47] = net320;
 assign la_data_out[48] = net321;
 assign la_data_out[49] = net322;
 assign la_data_out[4] = net277;
 assign la_data_out[50] = net323;
 assign la_data_out[51] = net324;
 assign la_data_out[52] = net325;
 assign la_data_out[53] = net326;
 assign la_data_out[54] = net327;
 assign la_data_out[55] = net328;
 assign la_data_out[56] = net329;
 assign la_data_out[57] = net330;
 assign la_data_out[58] = net331;
 assign la_data_out[59] = net332;
 assign la_data_out[5] = net278;
 assign la_data_out[60] = net333;
 assign la_data_out[61] = net334;
 assign la_data_out[62] = net335;
 assign la_data_out[63] = net336;
 assign la_data_out[6] = net279;
 assign la_data_out[7] = net280;
 assign la_data_out[8] = net281;
 assign la_data_out[9] = net282;
 assign user_irq[0] = net337;
 assign user_irq[1] = net338;
 assign user_irq[2] = net339;
 assign wbs_ack_o = net340;
 assign wbs_dat_o[0] = net341;
 assign wbs_dat_o[10] = net351;
 assign wbs_dat_o[11] = net352;
 assign wbs_dat_o[12] = net353;
 assign wbs_dat_o[13] = net354;
 assign wbs_dat_o[14] = net355;
 assign wbs_dat_o[15] = net356;
 assign wbs_dat_o[16] = net357;
 assign wbs_dat_o[17] = net358;
 assign wbs_dat_o[18] = net359;
 assign wbs_dat_o[19] = net360;
 assign wbs_dat_o[1] = net342;
 assign wbs_dat_o[20] = net361;
 assign wbs_dat_o[21] = net362;
 assign wbs_dat_o[22] = net363;
 assign wbs_dat_o[23] = net364;
 assign wbs_dat_o[24] = net365;
 assign wbs_dat_o[25] = net366;
 assign wbs_dat_o[26] = net367;
 assign wbs_dat_o[27] = net368;
 assign wbs_dat_o[28] = net369;
 assign wbs_dat_o[29] = net370;
 assign wbs_dat_o[2] = net343;
 assign wbs_dat_o[30] = net371;
 assign wbs_dat_o[31] = net372;
 assign wbs_dat_o[3] = net344;
 assign wbs_dat_o[4] = net345;
 assign wbs_dat_o[5] = net346;
 assign wbs_dat_o[6] = net347;
 assign wbs_dat_o[7] = net348;
 assign wbs_dat_o[8] = net349;
 assign wbs_dat_o[9] = net350;
endmodule

